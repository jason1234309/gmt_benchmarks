module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AMUX;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5Q;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5Q;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5Q;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CLK;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CLK;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D5Q;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CLK;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CLK;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AMUX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BMUX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CLK;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CLK;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CLK;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CLK;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CLK;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CLK;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B5Q;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A5Q;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B5Q;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BMUX;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5Q;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5Q;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CE;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_SR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BMUX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CLK;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CMUX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CLK;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AMUX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CE;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CLK;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_DO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_SR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CLK;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_DO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CLK;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D5Q;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DMUX;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BMUX;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CLK;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_DO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CLK;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CLK;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_DO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_AO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_AO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_AQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_BO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_BO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_CLK;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_CO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_CO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_CQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_DO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_DO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A5Q;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AMUX;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AX;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_BO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_BO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_BQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_CLK;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_CO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_CO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_CQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_DO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CLK;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BMUX;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CLK;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DMUX;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A5Q;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CLK;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CLK;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CLK;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AMUX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BMUX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CE;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CLK;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CMUX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_SR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CLK;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AMUX;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CLK;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_DO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CLK;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CLK;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CLK;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BMUX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CLK;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AMUX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BMUX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CE;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CLK;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DMUX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_SR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CLK;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CLK;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AMUX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BMUX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CLK;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CLK;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CLK;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C5Q;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A5Q;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CLK;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CLK;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DMUX;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D5Q;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A5Q;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C5Q;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A5Q;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A5Q;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AMUX;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AMUX;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AMUX;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AMUX;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CLK;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CLK;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CLK;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CLK;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B5Q;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B5Q;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CMUX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B5Q;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BMUX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B5Q;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CLK;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CLK;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AMUX;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AX;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BMUX;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CLK;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C5Q;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D5Q;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A5Q;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C5Q;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CE;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_SR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_AO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_AO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_BMUX;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_BO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_BO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_CLK;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_CO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_CO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_DO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_DO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_AO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_AO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_BO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_BO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_CO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_CO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_DO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_DO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AMUX;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_DO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_AO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_AO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_AQ;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_BO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_BO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_BQ;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_CLK;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_CO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_CO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_CQ;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_DO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_DO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_BO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_BO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_BQ;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CLK;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CQ;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_DO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_DO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_DQ;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_AO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_AO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_AQ;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_BO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_BO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_CLK;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_CO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_CO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_DO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_DO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A5Q;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AMUX;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AX;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_BMUX;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_BO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CLK;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_DO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_AO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_AO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_AQ;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_BO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_BO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_BQ;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_CLK;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_CO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_CO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_DO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_DO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_BO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CLK;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CMUX;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_DMUX;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A5Q;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AMUX;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AQ;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AX;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_BMUX;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_BO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CLK;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_DO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_BO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_BO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CLK;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CQ;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_DO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_DQ;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_AO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_AO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_BO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_BO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_CO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_CO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_DO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CLK;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_DO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_BO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CLK;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_DO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CLK;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_DO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CLK;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_DO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_BO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_DO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_AO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_AO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_BO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_BO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CMUX;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_DO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_DO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BMUX;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CLK;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CMUX;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_DMUX;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_DO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_BMUX;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_BO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CLK;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_DO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_DO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AMUX;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BMUX;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DMUX;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CLK;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_DO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CLK;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CLK;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_DO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D_XOR;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_A;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_A1;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_A2;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_A3;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_A4;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_A5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_A6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_AMUX;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_AO5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_AO6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_A_CY;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_A_XOR;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_B;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_B1;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_B2;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_B3;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_B4;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_B5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_B6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_BO5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_BO6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_B_CY;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_B_XOR;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_C;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_C1;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_C2;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_C3;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_C4;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_C5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_C6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_CO5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_CO6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_C_CY;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_C_XOR;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_D;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_D1;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_D2;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_D3;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_D4;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_D5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_D6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_DO5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_DO6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_D_CY;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X36Y143_D_XOR;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_A;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_A1;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_A2;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_A3;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_A4;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_A5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_A6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_AO5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_AO6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_A_CY;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_A_XOR;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_B;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_B1;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_B2;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_B3;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_B4;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_B5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_B6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_BO5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_BO6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_B_CY;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_B_XOR;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_C;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_C1;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_C2;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_C3;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_C4;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_C5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_C6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_CO5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_CO6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_C_CY;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_C_XOR;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_D;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_D1;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_D2;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_D3;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_D4;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_D5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_D6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_DO5;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_DO6;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_D_CY;
  wire [0:0] CLBLM_R_X25Y143_SLICE_X37Y143_D_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_AO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_BO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_BO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_CO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_CO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_DO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_DO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_AO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_AO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_BO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_BO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_CO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_CO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_DO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_DO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5Q;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CLK;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CLK;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5Q;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CLK;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CLK;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AMUX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AMUX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DMUX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A5Q;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A5Q;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AMUX;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B5Q;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BMUX;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BMUX;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AMUX;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CLK;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CMUX;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A5Q;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5Q;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B5Q;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BMUX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B5Q;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BMUX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5Q;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DMUX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa22222222)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffdffffffdd)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeefffffffcff)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_ALUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefffffffcffff)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_ALUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffffffffffddff)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaff000030303030)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_C5Q),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_A5Q),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc0c088bb88bb)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_DO6),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffe000ee00e0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00faf0faf0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0313000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_C5Q),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f00aaaacccc)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafeaa00005400)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I2(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddd88d8d8d888)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff77333733)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_C5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_A5Q),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaac3cc0000)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_CQ),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_DO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdd880000dd88)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_BLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffc00fc00fc00)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_D5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_BO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffbbffffffffff)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_DLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_CQ),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9f00900fcf00c00)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_BLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_DO6),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_CQ),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddddcc00111100)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO5),
.I4(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_A5Q),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h006a00aa00aa00aa)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I5(CLBLM_L_X12Y117_SLICE_X17Y117_CO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ffffaa00)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_CO6),
.I2(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_CQ),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3aca0a0acaca0a0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'habba0330f000f000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X17Y117_CO6),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X9Y119_BO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_DO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888dd88d8d8d8d8)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_DQ),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1b1b1a0a0a0a0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f044f044)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_CQ),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaff5000fa0050)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I1(1'b1),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_DQ),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_DO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcceeccec00220020)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_CQ),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000ffee5544)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_CQ),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0ffa0a0c0c0c0c0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_D5Q),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88b888bb88b888)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff88ff8800880088)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_DQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff144400001444)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_B5Q),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffececa0a0a0a0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_DQ),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cac0aa00aa00)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_AO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_BO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf011f011f011f011)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_D5Q),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8ffa8a8a8a8a8)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0c0f0c0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffc00fc00fc)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_AO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_CO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_DO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fc0ccacacaca)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2c0c0c0c0c0c0c0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_B5Q),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaafeaa44005400)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I2(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88b888bb88b888)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_CO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffffefff)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd8ffd800d800d8)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_CQ),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd888888888888888)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_A5Q),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0ccf0cc)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fdf55dd0fcf00cc)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_DLUT (
.I0(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_DQ),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_B5Q),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffae)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_CLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_AO6),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_AO6),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_DO6),
.I5(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h111f000f11110000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_BLUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I2(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I2(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdc)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_DLUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I3(CLBLL_L_X4Y123_SLICE_X4Y123_CO6),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_CO6),
.I5(CLBLL_L_X4Y123_SLICE_X4Y123_BO6),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000cc505050dc)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_CLUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I4(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I5(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000303055007530)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_BLUT (
.I0(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I1(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I5(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaeaaae000caaae)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_A5Q),
.I1(LIOB33_X0Y67_IOB_X0Y68_I),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33bb00aa33bb00aa)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_AO5),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010111110100000)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_CLUT (
.I0(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_BLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.I1(CLBLL_L_X4Y123_SLICE_X4Y123_DO6),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I3(CLBLM_R_X3Y123_SLICE_X2Y123_CO6),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_DO5),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_CO6),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h040404040404ff04)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_ALUT (
.I0(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I5(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000005000c0c0d0c)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_DLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_A5Q),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff3bff0a)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.I3(CLBLL_L_X4Y123_SLICE_X4Y123_AO6),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I5(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000004000)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7ffffffffef)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_AO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_BO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500050037330500)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_DLUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I5(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002030200)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcc0100cecc0200)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fffc00fc)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_BQ),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff22ff22fff2fff2)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_DLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004400000050)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_CQ),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefffefeeeeffee)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_BLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_DO6),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_AO6),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_AO6),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000430fffffeff)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f0f0fff5fff0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_DLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_AO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_DO6),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5d5d5dff0c0c0c)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_CLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_AO6),
.I1(LIOB33_X0Y63_IOB_X0Y63_I),
.I2(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.I3(CLBLM_R_X25Y143_SLICE_X36Y143_AO6),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_DQ),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000080000)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_AO6),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_AO6),
.I4(CLBLM_R_X5Y122_SLICE_X7Y122_CO6),
.I5(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_DLUT (
.I0(CLBLM_R_X3Y125_SLICE_X2Y125_DO6),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_CO6),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_CO5),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_DO6),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff1f0f11001100)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(LIOB33_X0Y67_IOB_X0Y67_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffff00980000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeffffffff7ffff)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004000000)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_DLUT (
.I0(CLBLM_R_X3Y125_SLICE_X2Y125_DO6),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_CO6),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_CO6),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_DO5),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffbffffff)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_CLUT (
.I0(CLBLM_R_X3Y125_SLICE_X2Y125_DO6),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_CO6),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_CO6),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfbbffffafaa)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_BLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_CO6),
.I1(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_AO6),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_DO6),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_ALUT (
.I0(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_CO5),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_BO6),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_DO5),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_DO6),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_CO6),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_AO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_BO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bb8bb88bb88bb88)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_BLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff28ffa02828a0a0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I5(CLBLM_R_X5Y122_SLICE_X6Y122_A5Q),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_AO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfffdff00008080)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffeff00004100)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbffffffffffbf)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_BLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff040004ff400040)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_C5Q),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888b8b8b8b8)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_ALUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff331100003311)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_CQ),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050005)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaa55001100)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_CLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33dd11cc00cc00)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc00cc50cc00)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f00aaaa0c00)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_DQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_DQ),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a0a3a0a3a3a3a3)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffe040000fe04)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafe005403030303)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_DQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I4(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_DO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3300aaaa3000)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_DLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5f0fa0005000a)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_CLUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacac0aaaaaa00)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaeeea55504440)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5fff5c00000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_DLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_CO6),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_DO6),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5f5a0a0a0a0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22fe32ee22ce02)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_BQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_CO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_AO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_BO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2442244242244224)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_CQ),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcac0cac00000aaaa)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_A5Q),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffe0ef000f404)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfff0aaa0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_CO6),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_AO6),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_BO6),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc08fc0000000000)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I3(CLBLM_L_X8Y118_SLICE_X11Y118_DO6),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha857a85703030303)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_CLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_CO6),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d888d8d888d88)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_A5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_DO6),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'habab0101baba1010)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_CO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_BO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_CO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fffdf5f5)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_CO5),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_B5Q),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffc00000f0c)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_DQ),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffccf0c0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_BLUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_DO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa003300cc)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_ALUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_BO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc00fc0000ff55ff)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_DQ),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f0fcccc0f00)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_CQ),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_CQ),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888dd88dd8888)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddd88d8d8d888)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_BO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_CO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf909fa0afa0afa0a)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_DLUT (
.I0(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a3a0a3a3a0a3a0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_CLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000eeee4444)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddd8d8dd88d888)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_BO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_CO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc0c0ffffcfc0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fef0fe000e000e)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_CLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_CQ),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00bb11aa00aa00)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_A5Q),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_BO6),
.I5(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff88ff8800880088)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_CO5),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_AO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_BO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_CO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_DO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fff0f03300)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_D5Q),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_B5Q),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f03300aaaaf0ff)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_CLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1a0e4a0b1a0e4)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaab0001aaaa0000)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I5(RIOB33_X105Y119_IOB_X1Y119_I),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_CO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeece00000050)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_DLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_DQ),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fef0fe000e000e)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_D5Q),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddcdc11111010)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_BLUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_DQ),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaffaaf0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_ALUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_BO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdffffff)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_DLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_CO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I3(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffd00aa00aa)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_CLUT (
.I0(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ee44ee44)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfecccc00320000)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_A5Q),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_BO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699669966996)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_DLUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e0f0a0a0a3a0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff660066ff000000)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfecc3200fecc3200)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_DO5),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_CO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_DO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5050f0f0ff00)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff9cff9c)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafc0cfc0c)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_BLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_DQ),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccf0cc00cc00)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_CO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a3a3acac)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_DLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafc00)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_CLUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a0e4f5e4a0e4)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_CQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffcec3020)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_DO6),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_BO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_CO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ccccf0f0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00cccc)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055ff44cc)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fc00fc00)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_BO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_CO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_DO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0030303030)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_DQ),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0f0c0f0c)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I1(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fff4fc050f040c)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I1(CLBLM_L_X8Y123_SLICE_X11Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbbbbbbbb8b)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_CO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_BO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_DO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfcfc00003030)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050cccccc00)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_B5Q),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0eef000f0ee)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaffaaf0aa00)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_ALUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_BO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000011001100)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeeaffff4440)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffff13333333)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_C5Q),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_CO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0aca3a0a0a3ac)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_CO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f011444444)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_BO5),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0e4e4f5a0e4e4)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaafe00540054)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_DQ),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_CO5),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_CO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acfc0cfc0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_CLUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8dd8f000f000)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1c0f3c0e2c0c0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.I4(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X10Y126_BO5),
.Q(CLBLM_L_X8Y126_SLICE_X10Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X10Y126_AO6),
.Q(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h337f337f7f7f7f7f)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_DLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_CLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h404000008888dd88)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_C5Q),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f88f888f888f888)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_AO5),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_AO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdddcfffa0000000)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_DO6),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I4(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888ff55aa00)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I4(RIOB33_X105Y125_IOB_X1Y126_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_BO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_CO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_DO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hceecceec0aa00aa0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_DLUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaccaacc)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_CLUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5b1b1b1a0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044faee5044)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaafbea11005140)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3ccc6ccc)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_BLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I5(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0ff05af0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I5(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_CO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555500000000)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_DLUT (
.I0(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc666ccccc)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I4(CLBLM_L_X8Y128_SLICE_X11Y128_DO6),
.I5(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc333633cc)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_BLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_AO5),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000110000005500)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_ALUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffcfcfc0c0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c4c444444444)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0054545454)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000fa00fa)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_ALUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_AO6),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f3f3c0c0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_C5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaa00cc)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddcdddc11101110)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_A5Q),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003322221111)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_DLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_C5Q),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h05fa00ff00ff00ff)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_CLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I3(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaaaaaa0000c000)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff400400004004)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffba008affba008a)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_CO5),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0023ff730023ff73)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_BO5),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h31000031ffceceff)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_C5Q),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_BO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_BO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_CO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_DO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafeaa00005400)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffc0e0d0f0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_CLUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_CO5),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I2(CLBLM_L_X12Y124_SLICE_X16Y124_BO6),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_DO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_AO6),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_DO6),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cc44cc44)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3336333355550000)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf10ef2010df20ef)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_AO6),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f470f8bf074f0b8)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_AO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_D5Q),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000330f000033a5)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_CQ),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555655ff33ff33)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_DQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_AO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_CO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa30aa30aa30aa30)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_DLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00d5d58080)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.I4(CLBLM_R_X13Y119_SLICE_X19Y119_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000e0e0e0e)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_BLUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000fcfc)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_AO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777bbbbddddeeee)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.I5(CLBLM_L_X12Y119_SLICE_X17Y119_A5Q),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff77bbffffddee)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_CLUT (
.I0(CLBLM_L_X12Y119_SLICE_X17Y119_BQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_C5Q),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_DQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h666606f66666f606)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_BLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_DQ),
.I1(CLBLM_L_X12Y119_SLICE_X17Y119_A5Q),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_AO6),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa0cc0000a0cc)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_CQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa20000aaaa0a0a)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0e000eff0f000f)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_CLUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_CO5),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I5(CLBLM_R_X13Y117_SLICE_X18Y117_AO6),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa0caa0faa0c)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcd0101dcdc1010)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y119_SLICE_X19Y119_AQ),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3ff3f3cfcffcfc)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_D5Q),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_CLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_A5Q),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I5(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000eee0000f000f)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc0ffc000c000c0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_DO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcec3020ffee3322)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_BO6),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8fcf8fc080c080c)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00bf15ea40)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hea40ff55ea40aa00)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffefffe)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_DLUT (
.I0(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_CQ),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000082824141)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_CLUT (
.I0(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_DQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000900900000000)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_BLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.I3(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_CO6),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f000acacacac)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_DQ),
.I1(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfefe00003232)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afafa0a0acac)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa008d888d88)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_DQ),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01ab01ba10ba10)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_A5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffeffffffff)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_DO6),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_BO6),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77dd77ff228822aa)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I1(CLBLM_L_X12Y119_SLICE_X17Y119_BQ),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I4(CLBLM_L_X12Y118_SLICE_X16Y118_DQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005555ff005050)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I3(CLBLM_L_X12Y118_SLICE_X16Y118_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f0ccf0ccf0cc)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_DLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff555500005555)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaabbaa11001100)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888e4a0e4a0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffafffffffa)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_DQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc00fc00f600fc00)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_C5Q),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_DO6),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_B5Q),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_A5Q),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_BO6),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_B5Q),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefeeebababaaa)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefeffffffffff)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_DLUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_B5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333332)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_CLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_CQ),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_DO6),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969966969969696)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_BO5),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_CQ),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_CO6),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbabaaaaa10100000)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_C5Q),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0323fff50303ffff)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_DQ),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010ffef01000100)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaffc800fa00c8)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_ALUT (
.I0(CLBLM_L_X8Y119_SLICE_X11Y119_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_CO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_DO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcac0cac0cac0cac0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0c00aaaa0c00)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_CLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a0e4f5e4a0e4)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haacfaa00aacfaaff)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0c0f0c0f0c0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_DLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_B5Q),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f1f2f102010201)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1a0a0b1b1a0a0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_BO6),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000e0eee0ee)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f2f2f202020202)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_DLUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404cfcfc0c0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I4(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccf0003ccfc0030)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3e2c0c0ffaa0000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_ALUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_C5Q),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_BO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_CO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaacfff)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0f0f02222)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_CLUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_C5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_DQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffea40ffffea40)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I4(CLBLM_R_X11Y123_SLICE_X14Y123_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa33aa30aa30)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_ALUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_CO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_DO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffc0cfe0efc0c)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_CO6),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacaff0ff000)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_CLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeae5404feae5404)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafeaaaa50540000)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_CO5),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_DO5),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaff00cccc)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_DLUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_C5Q),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1d1c0c0ffcc3300)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I4(CLBLM_R_X11Y120_SLICE_X15Y120_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcc0300ee22ee22)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccaaf0ccf0cc)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_DQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.R(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0f0fffbf)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_C5Q),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf1130eecf5530aa)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_BLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55a054a0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_ALUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_DO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff505000005050)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_DLUT (
.I0(CLBLM_R_X13Y125_SLICE_X18Y125_BO6),
.I1(1'b1),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f0fff000)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_CLUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeae0404ffaa5500)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555ffbf5515)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_DQ),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_BO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff0dff00ff)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_DLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_C5Q),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_CO6),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_DQ),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0a0f0a0000a000a)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f3f3d1d1)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_BLUT (
.I0(CLBLM_L_X10Y126_SLICE_X12Y126_DO6),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_DO6),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc50ff5000)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X13Y126_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.Q(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f5f1f5f0f5f1f5f)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_DLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_CO5),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffa00008888)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_CLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0c0c00000c0c)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h84cca5ff00cc00ff)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_CO6),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_AO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_BO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_CO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_DO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f044f044)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_DLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I2(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc1100ddcc1100)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_CLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffcc00003300)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.I4(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00f0005a)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_AO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_BO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_CO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h99999999a9a9a9a9)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_DLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3e2e2e2e2)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_CLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff220022ff220022)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_BLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_DQ),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc50ff5000)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f000f000f)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y128_SLICE_X12Y128_AO5),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h83c38bcf4703f4f3)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_ALUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_C5Q),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_AO6),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ffffefef)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777fffff0000000)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_C5Q),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I2(RIOB33_X105Y141_IOB_X1Y141_I),
.I3(RIOB33_X105Y139_IOB_X1Y140_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y115_SLICE_X16Y115_AO6),
.Q(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202131313020213)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_AO5),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(CLBLM_L_X12Y115_SLICE_X16Y115_BO6),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0044014511551054)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_CLUT (
.I0(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffffcc9ccccc)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_BLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff500050ff550055)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_ALUT (
.I0(CLBLM_L_X12Y115_SLICE_X16Y115_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y115_SLICE_X17Y115_AO6),
.Q(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05ab01af05ab01)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_CO6),
.I3(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_DQ),
.Q(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.R(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_DO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_CO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cff3cffff3cff3c)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I3(CLBLM_L_X12Y119_SLICE_X16Y119_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_BO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200010303030)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_AO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X17Y116_AO6),
.Q(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X17Y116_BO6),
.Q(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X17Y116_CO6),
.Q(CLBLM_L_X12Y116_SLICE_X17Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa55554455)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_DLUT (
.I0(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.I1(CLBLM_R_X13Y117_SLICE_X18Y117_CO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y118_SLICE_X17Y118_CO6),
.I4(CLBLM_R_X13Y116_SLICE_X18Y116_CO6),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_DO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f3c0d1c0f3c0d1)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_CLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y117_SLICE_X19Y117_BQ),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_DO6),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_CO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f606f000f000)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_BLUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_AO5),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_BO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccceeec00002220)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_AO6),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_AO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_DO5),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_AO6),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_CO6),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_DO6),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f3f3c0c0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I3(CLBLM_R_X13Y118_SLICE_X18Y118_BQ),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_DO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf80d08f5f00500)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_BQ),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_CO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf0fafa0c000a0a)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_BLUT (
.I0(CLBLM_R_X13Y118_SLICE_X18Y118_DQ),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_BO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888dddd8888d8d8)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_BQ),
.I2(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_CQ),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_AO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X17Y117_AO6),
.Q(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00cccccccc)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_DLUT (
.I0(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.I4(CLBLM_R_X13Y116_SLICE_X18Y116_BO6),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_DO5),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_DO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa8aa800000000)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_R_X13Y117_SLICE_X18Y117_BO6),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_DO6),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I4(CLBLM_L_X12Y117_SLICE_X17Y117_BO5),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_DO5),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_CO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f0effeeffe)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_BLUT (
.I0(CLBLM_R_X13Y117_SLICE_X18Y117_DO6),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_BO6),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_BO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafafaffaaeaea)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_B5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_AO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y118_SLICE_X16Y118_AO6),
.Q(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y118_SLICE_X16Y118_BO6),
.Q(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y118_SLICE_X16Y118_CO6),
.Q(CLBLM_L_X12Y118_SLICE_X16Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y118_SLICE_X16Y118_DO6),
.Q(CLBLM_L_X12Y118_SLICE_X16Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00fe54fe54)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y119_SLICE_X17Y119_BQ),
.I2(CLBLM_L_X12Y118_SLICE_X16Y118_DQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_DO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaafe00540054)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y118_SLICE_X16Y118_CQ),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_CO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f4f405050404)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_BLUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I1(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_BO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000054545454)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I1(CLBLM_L_X12Y118_SLICE_X16Y118_DQ),
.I2(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_AO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y118_SLICE_X17Y118_AO6),
.Q(CLBLM_L_X12Y118_SLICE_X17Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y118_SLICE_X17Y118_BO6),
.Q(CLBLM_L_X12Y118_SLICE_X17Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0e0e0e0e0e0e0e)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_DLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_CQ),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_DO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_CLUT (
.I0(CLBLM_R_X13Y118_SLICE_X18Y118_BQ),
.I1(CLBLM_R_X13Y117_SLICE_X19Y117_BQ),
.I2(CLBLM_R_X13Y118_SLICE_X18Y118_DQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I4(CLBLM_L_X12Y118_SLICE_X17Y118_AQ),
.I5(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_CO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcf0f00c0c0000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_BO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaac0c0ff00)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y118_SLICE_X17Y118_AQ),
.I3(CLBLM_R_X13Y118_SLICE_X18Y118_BQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_AO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X16Y119_AO6),
.Q(CLBLM_L_X12Y119_SLICE_X16Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X16Y119_BO6),
.Q(CLBLM_L_X12Y119_SLICE_X16Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X16Y119_CO6),
.Q(CLBLM_L_X12Y119_SLICE_X16Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X16Y119_DO6),
.Q(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff400040)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y119_SLICE_X16Y119_CQ),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_L_X10Y120_SLICE_X13Y120_BO6),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_DO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f00aaaa0c00)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_CLUT (
.I0(CLBLM_R_X13Y120_SLICE_X19Y120_AQ),
.I1(CLBLM_L_X12Y119_SLICE_X16Y119_CQ),
.I2(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_CO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffe0ef000f404)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X12Y119_SLICE_X16Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_DQ),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_BO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dc10dd11dc10)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y119_SLICE_X16Y119_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I4(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_AO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y120_SLICE_X18Y120_CO6),
.Q(CLBLM_L_X12Y119_SLICE_X17Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X17Y119_AO6),
.Q(CLBLM_L_X12Y119_SLICE_X17Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X17Y119_BO6),
.Q(CLBLM_L_X12Y119_SLICE_X17Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X17Y119_CO6),
.Q(CLBLM_L_X12Y119_SLICE_X17Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c3ccc3c3c3cc)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y119_SLICE_X17Y119_CQ),
.I2(CLBLM_R_X13Y121_SLICE_X18Y121_DQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_BO6),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_DO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f000f000)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X12Y118_SLICE_X17Y118_BQ),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_CO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0eff0e000e000e)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.I1(CLBLM_L_X12Y119_SLICE_X17Y119_BQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_BO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffc800c8)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_ALUT (
.I0(CLBLM_L_X12Y120_SLICE_X17Y120_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y119_SLICE_X17Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_AO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_BO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_CO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_DO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fc000000fc)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_DQ),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_DO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00eeee)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_CO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54ae04ae04)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I3(CLBLM_R_X13Y118_SLICE_X18Y118_DQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_DQ),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_BO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc400c4ffc000c0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I5(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_AO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X17Y120_AO6),
.Q(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.Q(CLBLM_L_X12Y120_SLICE_X17Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000088000000)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_DLUT (
.I0(CLBLM_L_X12Y119_SLICE_X17Y119_AQ),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I3(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_DO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafafcfcfcf0)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_CQ),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccc0ccc0ccc0)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_BLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_A5Q),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_BO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdedf5a5cccc0000)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_ALUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.I2(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y123_SLICE_X17Y123_AO5),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_AO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X16Y121_BO6),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00003300ffffffff)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaeeeeeaea)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_CQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc00fafa0000)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_BLUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_DQ),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_CQ),
.I2(CLBLM_L_X12Y120_SLICE_X17Y120_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000033303330)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X17Y121_AO6),
.Q(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X17Y121_BO6),
.Q(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X17Y121_CO6),
.Q(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000300010303030)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_DLUT (
.I0(CLBLM_L_X12Y119_SLICE_X17Y119_AQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I2(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I3(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I4(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfcfc00003030)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_DO6),
.I3(1'b1),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000baea1040)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y121_SLICE_X17Y121_DO5),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000decc1200)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X17Y121_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X16Y122_AO6),
.Q(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X16Y122_BO6),
.Q(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X16Y122_CO6),
.Q(CLBLM_L_X12Y122_SLICE_X16Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X16Y122_DO6),
.Q(CLBLM_L_X12Y122_SLICE_X16Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafae0504aaaa0000)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_DO6),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X12Y122_SLICE_X16Y122_DQ),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5e4e4e4e4)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_BO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffe0ef000f404)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5cca0ccf5cca0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_DQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y122_SLICE_X15Y122_DQ),
.Q(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.R(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaafffeabffaa)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_DLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.I2(CLBLM_L_X12Y123_SLICE_X17Y123_DO6),
.I3(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.I4(CLBLM_R_X11Y122_SLICE_X15Y122_CQ),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00cc00fa00fa)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_CLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_CQ),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0c0f0c0f0f0a0a)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_DQ),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I3(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc50ff5000)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I1(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.I4(CLBLM_R_X11Y122_SLICE_X15Y122_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_BO6),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_CO6),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_DO6),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0faf00a000a00)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_DLUT (
.I0(CLBLM_R_X13Y119_SLICE_X19Y119_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_DO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000044444444)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_CO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaccaaf0aaf0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_BLUT (
.I0(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I5(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_BO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bbb8bb8888b888)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_ALUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_CQ),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_AO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X17Y123_AO6),
.Q(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X17Y123_BO6),
.Q(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.Q(CLBLM_L_X12Y123_SLICE_X17Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffe7fffffff)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_DLUT (
.I0(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I2(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I4(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_AO5),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_DO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafaeae05050404)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y124_SLICE_X17Y124_CO6),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I3(1'b1),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.I5(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_CO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888bbbb8888bb88)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_BLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_CO6),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I5(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_BO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aacc000f0000)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_DQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_AO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_AO6),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3131313131313131)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_BLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555bbba1110)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.I2(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I3(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I5(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X17Y124_AO6),
.Q(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X17Y124_BO6),
.Q(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000100000000)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_DLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.I2(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y124_SLICE_X19Y124_CO6),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc336633c6)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_CLUT (
.I0(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_CQ),
.I2(CLBLM_R_X13Y124_SLICE_X18Y124_DO6),
.I3(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.I4(CLBLM_L_X12Y124_SLICE_X17Y124_DO6),
.I5(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faaccaa00aacc)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_BLUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.I5(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff5000550050)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I1(1'b1),
.I2(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I5(CLBLM_L_X12Y118_SLICE_X17Y118_AQ),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_DO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4a4a4a4a0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_CQ),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_DO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0e4e4e4f5)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_CO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f033f0ee)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_AO5),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_AO6),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_BO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0f0a0f8acf8acf)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y125_SLICE_X15Y125_DO6),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_AO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X17Y125_AO6),
.Q(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2fdf758a23df758a)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_DLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_DO6),
.I4(CLBLM_L_X12Y125_SLICE_X17Y125_BO5),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_DO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff8cffcccc8c8c)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_CLUT (
.I0(CLBLM_R_X13Y125_SLICE_X18Y125_BO6),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_DQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I4(CLBLM_L_X12Y125_SLICE_X17Y125_DO6),
.I5(CLBLM_L_X12Y125_SLICE_X17Y125_BO6),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_CO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000cc11115555)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_BO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff0fccccf000)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y125_SLICE_X17Y125_CO6),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_AO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_C5Q),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.R(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.R(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2033200000330000)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_CLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_BO5),
.I3(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_CO6),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa0101e341e2e2)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000200)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_DO5),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_AO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88b8888b88b888b8)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_DLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.I5(CLBLM_R_X13Y125_SLICE_X19Y125_BO6),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa000033c3)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_CO6),
.I3(CLBLM_R_X13Y126_SLICE_X18Y126_BO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55fb51aa00)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_BO6),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_BO6),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccffccf0ccf0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_AO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c0c4c0c5f0f5f0f)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_ALUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_CO6),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_A5Q),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_BO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_AO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0f0fff0ff)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ccf5f5f5f5)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff8ff88f8f88888)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I1(LIOB33_X0Y51_IOB_X0Y51_I),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffea0000ffc00000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_ALUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_C5Q),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddfffffffcffff)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_DO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.Q(CLBLM_R_X3Y118_SLICE_X3Y118_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.Q(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.Q(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88000000a8a0a0a0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ebc3ebc3)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_DO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddcccccdddcdddc)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_DO6),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_CO6),
.I4(CLBLM_R_X5Y117_SLICE_X6Y117_DO6),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2a2f3f3a2a2f3f3)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_DO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa2200aaaaaaaa)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff20ff0020200000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h03a30faf0faf0faf)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_DO6),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5f57ffff5555)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddddddddffdf)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_A5Q),
.I4(LIOB33_X0Y53_IOB_X0Y53_I),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_A5Q),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31fd31cd01fd31)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I4(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_A5Q),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdecc1200decc1200)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_DO6),
.I4(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffff55005555)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.Q(CLBLM_R_X3Y120_SLICE_X3Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.Q(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777070769966996)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I4(CLBLM_R_X3Y125_SLICE_X3Y125_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d800f00000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f2030200aa00aa)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e2e2ff00aaaa)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.Q(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88ddd8d88888d8d8)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500454405000500)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_ALUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I3(LIOB33_X0Y71_IOB_X0Y71_I),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_CQ),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000a0a00000f00)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_DLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_CQ),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff22f2ffff22f2)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_CLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I2(LIOB33_X0Y57_IOB_X0Y57_I),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_AO6),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000022ffff0f0f)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_ALUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_DO6),
.I1(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I4(CLBLM_R_X3Y124_SLICE_X3Y124_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff22f222f2)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_CO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y123_SLICE_X2Y123_BO6),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000c202)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_DQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d5d0c0cff5dff0c)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_ALUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I3(LIOB33_X0Y55_IOB_X0Y55_I),
.I4(LIOB33_X0Y61_IOB_X0Y61_I),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbfafabbfbaafa)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_DLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_AO5),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_C5Q),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_CLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I1(CLBLM_R_X3Y123_SLICE_X2Y123_AO6),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_DO6),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_DO6),
.I4(CLBLM_R_X7Y123_SLICE_X9Y123_BO6),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_DO6),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a2008000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I5(CLBLM_R_X3Y124_SLICE_X3Y124_AO6),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdffffffefff)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h75ff757530ff3030)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_DLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_CO5),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.I2(LIOB33_X0Y59_IOB_X0Y59_I),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I4(LIOB33_X0Y69_IOB_X0Y70_I),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7ffffffff7)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ffffffccccffff)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbffffffffffffbf)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_ALUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffa)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_CLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_DO6),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_CO6),
.I4(CLBLM_R_X3Y124_SLICE_X3Y124_BO6),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_BO6),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff88f8)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.I1(CLBLM_R_X25Y143_SLICE_X36Y143_AO6),
.I2(LIOB33_X0Y53_IOB_X0Y54_I),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_DO6),
.I5(CLBLM_R_X3Y126_SLICE_X2Y126_CO6),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbfffff)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccfccffdddfddff)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_DLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I1(CLBLM_R_X25Y143_SLICE_X36Y143_AO6),
.I2(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h05000d0c00000c0c)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_CLUT (
.I0(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I1(LIOB33_X0Y69_IOB_X0Y70_I),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I4(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdccccccccccccc)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X25Y143_SLICE_X36Y143_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefffe)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_ALUT (
.I0(CLBLM_R_X3Y126_SLICE_X2Y126_BO6),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_BO6),
.I2(CLBLL_L_X4Y124_SLICE_X4Y124_DO6),
.I3(LIOB33_X0Y59_IOB_X0Y59_I),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.I5(CLBLM_R_X3Y125_SLICE_X2Y125_CO6),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033323332)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_DLUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_BO6),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_CO6),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_DO6),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffbffffff)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_CLUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_AO6),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_CO6),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_BLUT (
.I0(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_BO6),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_AO6),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_CO6),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000100)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_DO6),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_CO6),
.I2(CLBLM_R_X3Y125_SLICE_X2Y125_AO6),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_BO6),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_CO6),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_CO6),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffffffffff)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000004000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(CLBLM_R_X25Y143_SLICE_X36Y143_AO6),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4f4f4f4f4fff4)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_BLUT (
.I0(CLBLM_R_X3Y126_SLICE_X2Y126_DO6),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(CLBLM_R_X3Y126_SLICE_X2Y126_AO6),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbffffffffffbfb)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(1'b1),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0044000000470003)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_AO5),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.I4(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300030370300000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_CLUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbfb08080808)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a8a8a8affffcfcf)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(1'b1),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_DO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_CO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_BO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdfffffffd)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_AO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_DO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_CO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_BO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafffffffff5f5)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(1'b1),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(1'b1),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_AO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfff5f002a00aa)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f099f000f000)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01144f0f00000)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f03030)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf444f555f444f444)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca0f0a0f0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_BO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00022aa00aa00)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000006666)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_BLUT (
.I0(CLBLM_R_X7Y118_SLICE_X9Y118_BQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50fa50ee44)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X7Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00055ff55ff)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h313330330f0f0000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_CLUT (
.I0(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cc00aaf0aaf0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_BLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff51ff4151514141)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cfc0cfc0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff03ff0c0003000c)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_CO6),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffee0044)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e4e4cccc)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X7Y118_AO6),
.Q(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.Q(CLBLM_R_X5Y118_SLICE_X7Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfdfcfdf0f1f0f1)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_DO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_BO6),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f1f1f1fff0f0f0f)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaabbee00001144)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_CQ),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaa0aaa0aaa0)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.I4(CLBLM_L_X12Y118_SLICE_X17Y118_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_BO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h400040000fff0fff)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I3(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0012122222)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd888d888d8)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.Q(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.Q(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aafe0054)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_DO6),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f5f400000504)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_DO6),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaa0aaa0aaa0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_CO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888fa50fa50)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00aaf0aaf0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_CLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0033aaaa00cc)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_DO6),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeaeeeaccc0ccc0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50dcf0fcdcdcfcfc)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_DLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f30000f5ff0000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_CLUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_DO6),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_DO6),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffbffffff)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccf0ccf0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.I2(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_AO5),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_BO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_CO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_DO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fe32cc00dc10)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaa0caafcaa0c)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff005454fcfc)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aacc0fcc0f)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_ALUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbfffffffb)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_DLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_CO6),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_C5Q),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_A5Q),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_A5Q),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_A5Q),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_A5Q),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_A5Q),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_D5Q),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_AO5),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffee)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_ALUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_A5Q),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_A5Q),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_BO5),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_BO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_CO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_CO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_CO6),
.I2(CLBLL_L_X4Y122_SLICE_X5Y122_CO6),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_DO6),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeff4455eeaa4400)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I4(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I5(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50fafa5050)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(RIOB33_X105Y127_IOB_X1Y127_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccfff000f0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_ALUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_B5Q),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00220022002f0022)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5fdfffff0fc)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_DO6),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.I4(CLBLM_R_X5Y122_SLICE_X7Y122_DO6),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_BLUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033500050)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_ALUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I5(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haabbbabbaaaababa)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I2(LIOB33_X0Y65_IOB_X0Y66_I),
.I3(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff757575ff303030)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_CLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_D5Q),
.I4(CLBLM_R_X25Y143_SLICE_X36Y143_AO6),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h004400440f4f0044)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_BLUT (
.I0(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeffffffeff)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_AO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbaffffffbaba)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_CO6),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_CO6),
.I4(CLBLM_R_X5Y122_SLICE_X7Y122_BO6),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000a000c)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000335000000050)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88d8d8d8d8)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff50ffdc)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_DLUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I2(LIOB33_X0Y65_IOB_X0Y65_I),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_CO6),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_AO5),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_CO6),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffbfa)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_CLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_BO6),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_BO6),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_BO6),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111000011f100f0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_DO6),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000fffc3330)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_A5Q),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_AO5),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ccafef00cca0ec)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_DLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_C5Q),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffdfffc)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_CLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_DO6),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_DO6),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_DO6),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_DO6),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffcf00500030)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_BLUT (
.I0(CLBLM_R_X3Y126_SLICE_X2Y126_DO6),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaf0f0ff00)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_A5Q),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_AO5),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff2fff2f2)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_CO6),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_BO6),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_DO6),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_DO6),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf00cf008a8a8a8a)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_CLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aac0aaf0aac0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0affc0ffc0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff2)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_DLUT (
.I0(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_DO6),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_CO6),
.I4(CLBLL_L_X4Y125_SLICE_X4Y125_CO6),
.I5(CLBLM_R_X5Y122_SLICE_X7Y122_AO6),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002020300)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_CLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005d0c00005500)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_BLUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffcfffcf)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_BO6),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_AO6),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30ff3030baffbaba)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_CLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_CO6),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_AO5),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303000003ab00aa)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_DO6),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffe)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_BO6),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_CO6),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_DO6),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_CO6),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000054045404)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_DLUT (
.I0(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000300022)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055307500003030)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_DO6),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7fdfdfffff)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_CO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080808080808080)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_DLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ba10aa00ea40)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_DQ),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_DO6),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3a0eca0eca0eca0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0012120000)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_ALUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_BO5),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_CO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_DLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0004400004444)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_CLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a3aca0a0a0a0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_A5Q),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_BO6),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f606f000f000)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_DO6),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_BLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0caa000000)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_BO6),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff2)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff000a)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_DLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff00fffffffc)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0d000000ff)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_BLUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00300000fcfc)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb000c00ff000000)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_DLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03030000a0a0afa0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0acafacacacacac)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaafc00)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.I2(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555551110000)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c00040ccc0ccc0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f10201f2f10201)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_BLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01122f0f01122)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_B5Q),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fff7fff)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffafffffffff)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_CO6),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0c0e0c0f0c0c0c)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_BLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf00a00fcfffcff)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_BO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_CO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1a0b1a0b1a0b1a0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffaaf0f0cc88)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_CO6),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeaccc0eeeaccc0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_ALUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.Q(CLBLM_R_X7Y118_SLICE_X9Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff0300fc0003)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000008000000)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_CLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_CQ),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4f1f104040101)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_DO5),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f404f101f404)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_DLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_CQ),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_BQ),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88e4e4e4e4)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_A5Q),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f2f1f201020102)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc50ccfacc50)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X9Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000036333333)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_DLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_A5Q),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_BQ),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbfbfb50505050)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00f0c0f0c0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_BQ),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5050ff50)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y119_SLICE_X17Y119_AQ),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffc)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_A5Q),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_C5Q),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_CO6),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_D5Q),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_AO6),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0002ffffffff)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaffabffaa)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_BO6),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_C5Q),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00a0cccc0000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_D5Q),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_BO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880000000000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_CLUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_DO6),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_DQ),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_DO6),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0ff4f40404)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_CO6),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff54fffc005400fc)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_D5Q),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffaa00f000aa)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffee0044)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaaaaaf8f88888)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555545400005454)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h070707070f0f0f00)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ee22ee22)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00088f0f00088)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_BQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeeec2220)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_C5Q),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_CO6),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_BO5),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cff0c0caeffaeae)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I5(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404fe0ef404)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_CLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafaaafcfc0c0c)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fafaf0f0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_CO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00220022000f0000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_DLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I3(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafae0504afae0504)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_D5Q),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0f404f404)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0aaaaaa)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_A5Q),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_BO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_CO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888880cff0c0c)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AO5),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1a0a0fa50fa50)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaccf0f0aacc)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_BLUT (
.I0(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3c0aaaaff00)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_CQ),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f2f2f2f22222222)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_DLUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AO5),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000000)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I5(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55dd00ccf5fdf0fc)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_BLUT (
.I0(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h73735050ff73ff50)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_ALUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_BQ),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_CO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h54550000fcff0000)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0e4e4e4e4)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005454ff005454)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_BLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fa50fa50)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f0f0f33330000)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300bfafb3a0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_CLUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0acacacac)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_BLUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_C5Q),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf5a0ff00)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I3(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05ae04af05ae04)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_D5Q),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fcfc0f000c0c)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_A5Q),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d8d8d8d8888888d)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_A5Q),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_DO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0fff000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_DLUT (
.I0(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcaca0000caca)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_C5Q),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00c0aaaa00c0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_BLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaacccc)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f005000af005100)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_DLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300c400cc00cc00)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_CLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_C5Q),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fc33ccf0f00000)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_BO5),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaba30300000ff00)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_ALUT (
.I0(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_CO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa000000aa000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_DLUT (
.I0(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffee00005544)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_A5Q),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I5(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf666f666f000f000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_DO6),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdefc5af0cccc0000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_ALUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_BQ),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888ddd8888888d8)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h04040404000f0000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_DLUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fffd00020002)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_CLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303fc0cf000f000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_CO6),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf909fa0af000f000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_ALUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_CO6),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f0000)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040000)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_C5Q),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccafafccccfafa)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_CO6),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0b4f0ffffccff)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_BO6),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00cc00c9)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050511114411)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaaf3f3)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_BLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_B5Q),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y115_SLICE_X14Y115_CO6),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h555655550f0f0000)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_BO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111111150505050)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_D5Q),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaffffff00f708)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_CLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05500f0f05555)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_BLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf888ff88ff88f888)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I3(CLBLM_L_X12Y124_SLICE_X16Y124_BO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_AO6),
.I5(CLBLM_R_X11Y115_SLICE_X14Y115_DO6),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_BO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_CO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0101313101023132)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_DLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafaff00005055)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_DO6),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacf0faaaac000)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_BLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd1111dcdc1010)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X15Y116_BO6),
.Q(CLBLM_R_X11Y116_SLICE_X15Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000006500ff0065)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_DLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_CQ),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_DQ),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000f02020d0d)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_CLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_BQ),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_A5Q),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00bbbb)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y123_SLICE_X11Y123_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y116_SLICE_X15Y116_CO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f2d0f0f00550055)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_BO5),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_BO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heefceefceefceecc)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffccffaaffc0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_CLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hea40ea40dddd8888)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafff0ccc0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_AO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699669999669966)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_DLUT (
.I0(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y119_SLICE_X16Y119_BQ),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bde7bde7bde7bde)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_CLUT (
.I0(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.I2(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_CQ),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffe0ff00ffe0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_CQ),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_AO5),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_BO5),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_BO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_CO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000000000)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_DLUT (
.I0(CLBLM_R_X13Y119_SLICE_X19Y119_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeaff44ff40)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_CQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_D5Q),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0a0a0fcfc0c0c)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffaa00aa)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_ALUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_B5Q),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_L_X12Y119_SLICE_X16Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3f3c3f3c3c3c3c)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I2(CLBLM_L_X12Y119_SLICE_X16Y119_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_BO6),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I2(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AO5),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc00fd0000005500)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_BLUT (
.I0(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_DQ),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffa8000000a8)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X11Y118_SLICE_X14Y118_CQ),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff3333ffff)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafa)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X13Y121_SLICE_X18Y121_DQ),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_BLUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_DO6),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_DQ),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_DO6),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_CO6),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc00fafa0000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_DQ),
.I1(CLBLM_L_X12Y119_SLICE_X16Y119_BQ),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_AO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_DQ),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y119_SLICE_X17Y119_CQ),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0eef000f0ee)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_CLUT (
.I0(CLBLM_L_X12Y119_SLICE_X16Y119_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_B5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1a0b1a0bb11aa00)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_BQ),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_CQ),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_DQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbaba11111010)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_CQ),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_BO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0054545454)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_DO6),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_DQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaac0ccccc0c0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_CLUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddccee00110022)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_CO5),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dc10cc00cc00)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I3(CLBLM_L_X12Y119_SLICE_X16Y119_CQ),
.I4(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_BO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_CO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_DO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fc30cc00fc30)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_A5Q),
.I3(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fc30cc00fc30)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_DQ),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ff55aa00)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I3(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I4(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe00feff100010)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_CQ),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011001100000000)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff9ffffffffff)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_CLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_AO5),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_DO6),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_DO6),
.I5(CLBLM_L_X10Y121_SLICE_X13Y121_BO5),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000ccacacaca)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3e2c0c0ffaa0000)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_ALUT (
.I0(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y121_SLICE_X18Y121_DQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X15Y121_AO6),
.Q(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X15Y121_BO6),
.Q(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X15Y121_CO6),
.Q(CLBLM_R_X11Y121_SLICE_X15Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.Q(CLBLM_R_X11Y121_SLICE_X15Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fa50ee44ea40)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_DQ),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_DO6),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0e4a0a0a0a0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y121_SLICE_X15Y121_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_CQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_BQ),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000404ff00fefe)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y121_SLICE_X13Y121_BO6),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f000fff0a000a)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_ALUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_BO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_CO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f011221122)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_DLUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff11ff4400110044)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_DQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_BO5),
.I5(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54aa00fcfc0000)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000005a5a)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_ALUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.I3(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X15Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.Q(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X15Y122_CO6),
.Q(CLBLM_R_X11Y122_SLICE_X15Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X15Y122_DO6),
.Q(CLBLM_R_X11Y122_SLICE_X15Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00ccf0cc)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_DQ),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0aaf0ccf0aa)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_CLUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_CQ),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.I5(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0e4f0e4)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0022222020)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffcfffffffff)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_DQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff4fff4)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I2(CLBLM_L_X12Y123_SLICE_X17Y123_DO6),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_DO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_ALUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_DO6),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_BO6),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X15Y123_AO6),
.Q(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X15Y123_BO6),
.Q(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X15Y123_CO6),
.Q(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdffffffff)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_DLUT (
.I0(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0a0800000a08)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0cfc0cfc0c0)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00f0cccc)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_DQ),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_CO5),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_DO5),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_CO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_DO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_DLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I1(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_A5Q),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffffcc00)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_A5Q),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfc0030ccfc0030)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303f303f000f000)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_A5Q),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_CO5),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_DLUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44eeee4444)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y143_IOB_X1Y144_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000101ff006868)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_BLUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa30aa30aa03aa03)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X13Y120_SLICE_X19Y120_BO5),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_BO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55ea15aa55ea15)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_DLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_DO6),
.I3(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000031333122)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_CLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_C5Q),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0cff0c00)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00ccf0cc)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_DQ),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X15Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X15Y125_BO6),
.Q(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X15Y125_CO6),
.Q(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa5a595555)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_DLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_CO5),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_BO5),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d000d00dddddddd)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_DO6),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7700777733003333)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_BLUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_DO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaacca0cca0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X8Y126_SLICE_X10Y126_A5Q),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.R(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h444c000000002220)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00df00ff00f7)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_CLUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_CO6),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000002)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_BLUT (
.I0(CLBLM_L_X10Y126_SLICE_X12Y126_CO6),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500000400)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_ALUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_AO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3033333331333133)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_DLUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_CO5),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_BO5),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000003030)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_CLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_BO5),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088008800)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_BLUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I3(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb7b700b733330033)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_DO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y121_SLICE_X15Y121_DQ),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_BO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c6c3c3c6c3c3c3)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_DLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I5(CLBLM_L_X10Y126_SLICE_X12Y126_CO6),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00fe0000f1f1)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f3f3f300f300f3)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_DO6),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0bbb0bbb00bb00bb)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_ALUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_DO6),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X15Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa99aa55aa95)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_DLUT (
.I0(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_BO5),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a9a9a5a5a9a5)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_CLUT (
.I0(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_CO6),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_BO6),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000bbfb0000bfff)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_BLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I1(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_BO5),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb33bb33b0000b33b)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_ALUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I3(CLBLM_R_X11Y127_SLICE_X15Y127_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y116_SLICE_X18Y116_AO6),
.Q(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X18Y116_DO5),
.O6(CLBLM_R_X13Y116_SLICE_X18Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffccffcc)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.O5(CLBLM_R_X13Y116_SLICE_X18Y116_CO5),
.O6(CLBLM_R_X13Y116_SLICE_X18Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0e0f0f)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_BLUT (
.I0(CLBLM_R_X13Y117_SLICE_X18Y117_CO6),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I2(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I4(CLBLM_L_X12Y118_SLICE_X17Y118_CO6),
.I5(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.O5(CLBLM_R_X13Y116_SLICE_X18Y116_BO5),
.O6(CLBLM_R_X13Y116_SLICE_X18Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8bb888888bb88)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_ALUT (
.I0(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y116_SLICE_X18Y116_AO5),
.O6(CLBLM_R_X13Y116_SLICE_X18Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X19Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X19Y116_DO5),
.O6(CLBLM_R_X13Y116_SLICE_X19Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X19Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X19Y116_CO5),
.O6(CLBLM_R_X13Y116_SLICE_X19Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X19Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X19Y116_BO5),
.O6(CLBLM_R_X13Y116_SLICE_X19Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X19Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X19Y116_AO5),
.O6(CLBLM_R_X13Y116_SLICE_X19Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b7b7b7bdededede)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_DLUT (
.I0(CLBLM_R_X13Y119_SLICE_X19Y119_AQ),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_DO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefefffffefe)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_CLUT (
.I0(CLBLM_R_X13Y119_SLICE_X19Y119_AQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I2(CLBLM_L_X12Y117_SLICE_X16Y117_BQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y118_SLICE_X18Y118_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_CO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff5affff5a)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_BLUT (
.I0(CLBLM_R_X13Y118_SLICE_X18Y118_CQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I3(CLBLM_R_X13Y118_SLICE_X18Y118_DQ),
.I4(CLBLM_R_X13Y117_SLICE_X19Y117_AQ),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_CO6),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699669969669)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_BO6),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I4(CLBLM_R_X13Y117_SLICE_X19Y117_AQ),
.I5(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_AO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y117_SLICE_X19Y117_AO6),
.Q(CLBLM_R_X13Y117_SLICE_X19Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y117_SLICE_X19Y117_BO6),
.Q(CLBLM_R_X13Y117_SLICE_X19Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y117_SLICE_X19Y117_CO6),
.Q(CLBLM_R_X13Y117_SLICE_X19Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_DO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaa00c0)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_CLUT (
.I0(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y117_SLICE_X19Y117_CQ),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_CO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccaaf0f000aa)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I1(CLBLM_R_X13Y117_SLICE_X19Y117_BQ),
.I2(CLBLM_R_X13Y117_SLICE_X19Y117_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_BO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300fedc3210)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y117_SLICE_X19Y117_AQ),
.I3(CLBLM_R_X13Y117_SLICE_X19Y117_CQ),
.I4(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_AO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y118_SLICE_X18Y118_AO6),
.Q(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y118_SLICE_X18Y118_BO6),
.Q(CLBLM_R_X13Y118_SLICE_X18Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y118_SLICE_X18Y118_CO6),
.Q(CLBLM_R_X13Y118_SLICE_X18Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y118_SLICE_X18Y118_DO6),
.Q(CLBLM_R_X13Y118_SLICE_X18Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000e444e444)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.I2(CLBLM_R_X13Y118_SLICE_X18Y118_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_DO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00c0c0aaaa)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_CLUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I1(CLBLM_R_X13Y118_SLICE_X18Y118_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_CO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f5a0a0a0f5a0)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y118_SLICE_X18Y118_BQ),
.I2(CLBLM_R_X13Y122_SLICE_X18Y122_CQ),
.I3(CLBLM_R_X13Y117_SLICE_X19Y117_BQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_BO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb100b1ff110011)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_ALUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_DO6),
.I2(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y118_SLICE_X19Y118_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_AO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y118_SLICE_X19Y118_AO6),
.Q(CLBLM_R_X13Y118_SLICE_X19Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_DO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_CO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_BO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fffc00f000fc)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X13Y118_SLICE_X19Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_AO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y119_SLICE_X18Y119_BO6),
.Q(CLBLM_R_X13Y119_SLICE_X18Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y119_SLICE_X18Y119_AO6),
.Q(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y119_SLICE_X18Y119_CO6),
.Q(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_DQ),
.I3(CLBLM_L_X12Y118_SLICE_X17Y118_BQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y119_SLICE_X19Y119_BQ),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_DO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00011f0f06688)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_CLUT (
.I0(CLBLM_L_X12Y118_SLICE_X17Y118_BQ),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_C5Q),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_CO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ddf0ee0000aaaa)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000120012)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_ALUT (
.I0(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_DO5),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_AO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y119_SLICE_X19Y119_AO6),
.Q(CLBLM_R_X13Y119_SLICE_X19Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y119_SLICE_X19Y119_BO6),
.Q(CLBLM_R_X13Y119_SLICE_X19Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_DO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_CO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11cc00dd11cc00)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_BO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb888bbbbb8888888)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y119_SLICE_X19Y119_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(CLBLM_R_X13Y118_SLICE_X18Y118_CQ),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_AO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y120_SLICE_X18Y120_AO6),
.Q(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y120_SLICE_X18Y120_BO6),
.Q(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100010000000100)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_DLUT (
.I0(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_A5Q),
.I2(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I4(CLBLM_R_X13Y121_SLICE_X18Y121_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_DO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a011001100)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_CLUT (
.I0(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I4(CLBLM_R_X13Y120_SLICE_X19Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_CO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a3aca3ac)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_BLUT (
.I0(CLBLM_R_X13Y120_SLICE_X19Y120_A5Q),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_BO5),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_BO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ce02fc30)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_ALUT (
.I0(CLBLM_R_X13Y121_SLICE_X18Y121_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I3(CLBLM_R_X13Y117_SLICE_X19Y117_CQ),
.I4(CLBLM_R_X13Y120_SLICE_X18Y120_CO5),
.I5(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_AO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y120_SLICE_X19Y120_BO6),
.Q(CLBLM_R_X13Y120_SLICE_X19Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y120_SLICE_X19Y120_AO6),
.Q(CLBLM_R_X13Y120_SLICE_X19Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_DO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_CO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a8a857575757)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I2(CLBLM_R_X13Y120_SLICE_X19Y120_AQ),
.I3(CLBLM_R_X13Y118_SLICE_X18Y118_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_BO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccfff0ffccffa0)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I2(CLBLM_R_X13Y120_SLICE_X19Y120_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_AO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y121_SLICE_X18Y121_AO6),
.Q(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y121_SLICE_X18Y121_BO6),
.Q(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y121_SLICE_X18Y121_CO6),
.Q(CLBLM_R_X13Y121_SLICE_X18Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.Q(CLBLM_R_X13Y121_SLICE_X18Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00f0f0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_DO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaa33cc)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_CLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I1(CLBLM_R_X13Y121_SLICE_X18Y121_CQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_CO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf5f8f00d050800)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_BLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y118_SLICE_X17Y118_AQ),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_BO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafff0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_ALUT (
.I0(CLBLM_R_X13Y121_SLICE_X18Y121_CQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_AO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_DO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_CO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_BO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_AO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y122_SLICE_X18Y122_AO6),
.Q(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y122_SLICE_X18Y122_BO6),
.Q(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.Q(CLBLM_R_X13Y122_SLICE_X18Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff39ff3cff39ff3c)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_DLUT (
.I0(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.I1(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_DO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000ccf0f0aaaa)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_CLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I1(CLBLM_R_X13Y122_SLICE_X18Y122_CQ),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_CO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000cfafa0a0a)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_BLUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I1(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I4(CLBLM_R_X13Y119_SLICE_X19Y119_BQ),
.I5(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_BO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f2f2f202020202)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_ALUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_DO6),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_AO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y122_SLICE_X19Y122_AO6),
.Q(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_DLUT (
.I0(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_AO5),
.I2(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I4(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I5(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_DO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_CLUT (
.I0(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I2(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I3(CLBLM_R_X13Y126_SLICE_X18Y126_AO5),
.I4(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I5(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_CO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff10ff00ffd0)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_BLUT (
.I0(CLBLM_R_X13Y122_SLICE_X19Y122_DO6),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_DQ),
.I3(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.I5(CLBLM_R_X13Y122_SLICE_X19Y122_CO6),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_BO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ff55fa50fa50)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_AO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_AO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_BO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_DO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00d07f2f8)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_CLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_AO5),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I4(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I5(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_CO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0054545151)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_BLUT (
.I0(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cfcfff00dcdc)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_ALUT (
.I0(CLBLM_R_X13Y125_SLICE_X18Y125_DO6),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I2(CLBLM_R_X13Y120_SLICE_X18Y120_DO5),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_AO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X19Y123_AO6),
.Q(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X19Y123_BO6),
.Q(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X19Y123_CO6),
.Q(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haefbaffaaffaaffa)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_DLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I4(CLBLM_R_X13Y124_SLICE_X19Y124_BO6),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_DO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000b0bff000e0e)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_CLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.I1(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I3(CLBLM_L_X12Y123_SLICE_X16Y123_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y122_SLICE_X19Y122_BO6),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_CO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faf0fa000a000a)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_BLUT (
.I0(CLBLM_R_X13Y123_SLICE_X19Y123_DO6),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I4(1'b1),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_BO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8ddddd8d8d8d8)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_CQ),
.I2(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_AO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffffffffff)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_DLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I1(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.I2(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y124_SLICE_X18Y124_BO6),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_DO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_CLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I1(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.I2(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I4(CLBLM_L_X12Y123_SLICE_X17Y123_CQ),
.I5(CLBLM_R_X13Y124_SLICE_X18Y124_BO6),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_CO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808000008880000)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_BLUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I1(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_BO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000bbffbfbf)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_ALUT (
.I0(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I2(CLBLM_R_X13Y124_SLICE_X19Y124_CO6),
.I3(CLBLM_R_X13Y124_SLICE_X18Y124_BO6),
.I4(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_AO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_DO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004040400)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_CLUT (
.I0(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I2(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_CO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0000304c000020)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I4(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_BO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.I1(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.I2(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_CQ),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I5(CLBLM_R_X13Y124_SLICE_X19Y124_CO6),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_AO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y125_SLICE_X18Y125_AO6),
.Q(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h003300330f0f5f7f)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_DLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I2(CLBLM_R_X13Y120_SLICE_X18Y120_DO5),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_BO5),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7377777700880088)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_CLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I1(CLBLM_R_X13Y120_SLICE_X18Y120_DO5),
.I2(CLBLM_R_X13Y125_SLICE_X19Y125_BO5),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555000533333332)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I1(CLBLM_R_X13Y125_SLICE_X19Y125_BO5),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff541000005410)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X13Y125_SLICE_X19Y125_BO6),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_C5Q),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_AO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y125_SLICE_X19Y125_AO6),
.Q(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333c3cc3333c6cc)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_DLUT (
.I0(CLBLM_R_X13Y124_SLICE_X19Y124_AO6),
.I1(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.I3(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.I5(CLBLM_R_X13Y124_SLICE_X18Y124_CO6),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_DO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fff70000ffdf)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_CLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_CQ),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_AO5),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_CO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3330003033300030)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.I2(CLBLM_R_X13Y124_SLICE_X19Y124_AO6),
.I3(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_CO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_BO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f2f203030202)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_ALUT (
.I0(CLBLM_R_X13Y125_SLICE_X19Y125_DO6),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_AO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555455ffffffff)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_DLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I5(CLBLM_R_X13Y120_SLICE_X18Y120_DO5),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb773a55000000000)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_CLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_BO5),
.I5(CLBLM_R_X13Y125_SLICE_X19Y125_BO6),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_CO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000022220000)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I3(CLBLM_R_X13Y125_SLICE_X19Y125_BO6),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_BO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0dd0f0ff0f0f000)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_AO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X19Y126_AO6),
.Q(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_DO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_CO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_BO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbaab11111001)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I2(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I3(CLBLM_R_X13Y125_SLICE_X19Y125_CO6),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_AO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.Q(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff2aff28002a0028)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_CO6),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y130_SLICE_X18Y130_AO6),
.Q(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_DO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_CO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0ffaaaaf0f0)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_AO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_DO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_CO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_AO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y143_SLICE_X36Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y143_SLICE_X36Y143_DO5),
.O6(CLBLM_R_X25Y143_SLICE_X36Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y143_SLICE_X36Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y143_SLICE_X36Y143_CO5),
.O6(CLBLM_R_X25Y143_SLICE_X36Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y143_SLICE_X36Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y143_SLICE_X36Y143_BO5),
.O6(CLBLM_R_X25Y143_SLICE_X36Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbbffffffaa)
  ) CLBLM_R_X25Y143_SLICE_X36Y143_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(1'b1),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(1'b1),
.O5(CLBLM_R_X25Y143_SLICE_X36Y143_AO5),
.O6(CLBLM_R_X25Y143_SLICE_X36Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y143_SLICE_X37Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y143_SLICE_X37Y143_DO5),
.O6(CLBLM_R_X25Y143_SLICE_X37Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y143_SLICE_X37Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y143_SLICE_X37Y143_CO5),
.O6(CLBLM_R_X25Y143_SLICE_X37Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y143_SLICE_X37Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y143_SLICE_X37Y143_BO5),
.O6(CLBLM_R_X25Y143_SLICE_X37Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y143_SLICE_X37Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y143_SLICE_X37Y143_AO5),
.O6(CLBLM_R_X25Y143_SLICE_X37Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_DO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_CO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_BO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000a0a0a0a)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_ALUT (
.I0(RIOB33_X105Y119_IOB_X1Y119_I),
.I1(1'b1),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_AO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_DO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_CO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_BO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_AO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_ALUT (
.I0(RIOB33_X105Y139_IOB_X1Y139_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffaaaaffff)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffaaaaffff)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffff00ffff)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_ALUT (
.I0(CLBLM_R_X13Y118_SLICE_X19Y118_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffaaaaffff)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_L_X12Y117_SLICE_X16Y117_D5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_R_X7Y121_SLICE_X9Y121_CQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_L_X12Y117_SLICE_X16Y117_DQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_R_X5Y122_SLICE_X6Y122_B5Q),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X8Y126_SLICE_X11Y126_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X7Y121_SLICE_X9Y121_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X7Y122_SLICE_X8Y122_B5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_L_X10Y124_SLICE_X13Y124_D5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y118_SLICE_X3Y118_A5Q),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y138_SLICE_X163Y138_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_R_X11Y152_SLICE_X14Y152_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLM_R_X37Y120_SLICE_X56Y120_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_L_X12Y118_SLICE_X17Y118_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_BO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_CO6),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_CO5),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_R_X11Y152_SLICE_X14Y152_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X10Y130_BO6),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO6),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_L_X12Y130_SLICE_X16Y130_BO5),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_L_X12Y130_SLICE_X16Y130_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_L_X12Y118_SLICE_X17Y118_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_BO5),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_CO6),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_CO5),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X13Y118_SLICE_X19Y118_AQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X25Y143_SLICE_X36Y143_AO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X25Y143_SLICE_X36Y143_AO5),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_AMUX = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_AMUX = CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_BMUX = CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_AMUX = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D = CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D = CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_AMUX = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_CMUX = CLBLL_L_X4Y117_SLICE_X4Y117_C5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_DMUX = CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_CMUX = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_AMUX = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CMUX = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_AMUX = CLBLL_L_X4Y119_SLICE_X5Y119_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_AMUX = CLBLL_L_X4Y120_SLICE_X4Y120_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_BMUX = CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_AMUX = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A = CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A = CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_DMUX = CLBLL_L_X4Y121_SLICE_X5Y121_D5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_DMUX = CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A = CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A = CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B = CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C = CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_AMUX = CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_DMUX = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C = CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_AMUX = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_AMUX = CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A = CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B = CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C = CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A = CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C = CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_AMUX = CLBLL_L_X4Y125_SLICE_X4Y125_AO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A = CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_AMUX = CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_BMUX = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A = CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B = CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A = CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_BMUX = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_CMUX = CLBLL_L_X4Y127_SLICE_X5Y127_CO5;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_DMUX = CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_AMUX = CLBLM_L_X8Y115_SLICE_X11Y115_AO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_AMUX = CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_BMUX = CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_CMUX = CLBLM_L_X8Y116_SLICE_X11Y116_C5Q;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A = CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B = CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_AMUX = CLBLM_L_X8Y117_SLICE_X10Y117_A5Q;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_CMUX = CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_DMUX = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B = CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_CMUX = CLBLM_L_X8Y117_SLICE_X11Y117_CO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_DMUX = CLBLM_L_X8Y118_SLICE_X11Y118_DO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_DMUX = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A = CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B = CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C = CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A = CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_CMUX = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_DMUX = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C = CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_DMUX = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_CMUX = CLBLM_L_X8Y121_SLICE_X10Y121_CO5;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A = CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A = CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C = CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D = CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_DMUX = CLBLM_L_X8Y122_SLICE_X10Y122_D5Q;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A = CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B = CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A = CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A = CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A = CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B = CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C = CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_AMUX = CLBLM_L_X8Y124_SLICE_X10Y124_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_CMUX = CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A = CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A = CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B = CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A = CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B = CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_AMUX = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_BMUX = CLBLM_L_X8Y125_SLICE_X11Y125_BO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_CMUX = CLBLM_L_X8Y125_SLICE_X11Y125_C5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_AMUX = CLBLM_L_X8Y126_SLICE_X10Y126_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_BMUX = CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_DMUX = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A = CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B = CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_AMUX = CLBLM_L_X8Y126_SLICE_X11Y126_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_BMUX = CLBLM_L_X8Y126_SLICE_X11Y126_BO5;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A = CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B = CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C = CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D = CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A = CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B = CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A = CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B = CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C = CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D = CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A = CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B = CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C = CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_AMUX = CLBLM_L_X8Y128_SLICE_X11Y128_AO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A = CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C = CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_AMUX = CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_BMUX = CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_BMUX = CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B = CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C = CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D = CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_AMUX = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_AMUX = CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_CMUX = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A = CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B = CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A = CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A = CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_BMUX = CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_DMUX = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_AMUX = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_BMUX = CLBLM_L_X10Y119_SLICE_X12Y119_B5Q;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_CMUX = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_AMUX = CLBLM_L_X10Y120_SLICE_X12Y120_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_BMUX = CLBLM_L_X10Y120_SLICE_X12Y120_B5Q;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_CMUX = CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A = CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B = CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A = CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_BMUX = CLBLM_L_X10Y121_SLICE_X13Y121_BO5;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A = CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_AMUX = CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_DMUX = CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_AMUX = CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_CMUX = CLBLM_L_X10Y123_SLICE_X12Y123_C5Q;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_CMUX = CLBLM_L_X10Y123_SLICE_X13Y123_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A = CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B = CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CMUX = CLBLM_L_X10Y124_SLICE_X12Y124_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_AMUX = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_BMUX = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CMUX = CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_DMUX = CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A = CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_AMUX = CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A = CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A = CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_CMUX = CLBLM_L_X10Y126_SLICE_X12Y126_CO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A = CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_CMUX = CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_DMUX = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A = CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B = CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C = CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A = CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B = CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D = CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C = CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_AMUX = CLBLM_L_X10Y128_SLICE_X12Y128_AO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B = CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B = CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D = CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A = CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B = CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B = CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_AMUX = CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_BMUX = CLBLM_L_X12Y115_SLICE_X16Y115_BO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_CMUX = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A = CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B = CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C = CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A = CLBLM_L_X12Y116_SLICE_X16Y116_AO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B = CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D = CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_AMUX = CLBLM_L_X12Y116_SLICE_X16Y116_AO5;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A = CLBLM_L_X12Y116_SLICE_X17Y116_AO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B = CLBLM_L_X12Y116_SLICE_X17Y116_BO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C = CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D = CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C = CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D = CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_DMUX = CLBLM_L_X12Y117_SLICE_X16Y117_D5Q;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A = CLBLM_L_X12Y117_SLICE_X17Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B = CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D = CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_BMUX = CLBLM_L_X12Y117_SLICE_X17Y117_BO5;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A = CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C = CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D = CLBLM_L_X12Y118_SLICE_X16Y118_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A = CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B = CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C = CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A = CLBLM_L_X12Y119_SLICE_X16Y119_AO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B = CLBLM_L_X12Y119_SLICE_X16Y119_BO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C = CLBLM_L_X12Y119_SLICE_X16Y119_CO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D = CLBLM_L_X12Y119_SLICE_X16Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A = CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B = CLBLM_L_X12Y119_SLICE_X17Y119_BO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C = CLBLM_L_X12Y119_SLICE_X17Y119_CO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_AMUX = CLBLM_L_X12Y119_SLICE_X17Y119_A5Q;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A = CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B = CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C = CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D = CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A = CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_BMUX = CLBLM_L_X12Y120_SLICE_X17Y120_BO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_DMUX = CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_AMUX = CLBLM_L_X12Y121_SLICE_X16Y121_A5Q;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_BMUX = CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A = CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B = CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C = CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_DMUX = CLBLM_L_X12Y121_SLICE_X17Y121_DO5;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A = CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B = CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A = CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_AMUX = CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_BMUX = CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_CMUX = CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B = CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C = CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A = CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B = CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_AMUX = CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A = CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C = CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D = CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A = CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B = CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C = CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A = CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B = CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C = CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D = CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_BMUX = CLBLM_L_X12Y125_SLICE_X17Y125_BO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_AMUX = CLBLM_L_X12Y126_SLICE_X16Y126_AO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_BMUX = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_DMUX = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A = CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A = CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B = CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C = CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D = CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A = CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A = CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B = CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C = CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D = CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_AMUX = CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_BMUX = CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D = CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_AMUX = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_AMUX = CLBLM_R_X3Y118_SLICE_X3Y118_A5Q;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_CMUX = CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_AMUX = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_AMUX = CLBLM_R_X3Y120_SLICE_X3Y120_A5Q;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_BMUX = CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_CMUX = CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_DMUX = CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_AMUX = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_AMUX = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_AMUX = CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_DMUX = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_AMUX = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_BMUX = CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_CMUX = CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_AMUX = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_BMUX = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_CMUX = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A = CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_AMUX = CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_BMUX = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D = CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_AMUX = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_BMUX = CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B = CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C = CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D = CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_AMUX = CLBLM_R_X3Y127_SLICE_X3Y127_AO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_DMUX = CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_AMUX = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_CMUX = CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_BMUX = CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_CMUX = CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_DMUX = CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_CMUX = CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CMUX = CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_DMUX = CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CMUX = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_DMUX = CLBLM_R_X5Y120_SLICE_X6Y120_D5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A = CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_AMUX = CLBLM_R_X5Y121_SLICE_X6Y121_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_AMUX = CLBLM_R_X5Y121_SLICE_X7Y121_AO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A = CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B = CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_AMUX = CLBLM_R_X5Y122_SLICE_X6Y122_A5Q;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_BMUX = CLBLM_R_X5Y122_SLICE_X6Y122_B5Q;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A = CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B = CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_BMUX = CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B = CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C = CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_AMUX = CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A = CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B = CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C = CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_CMUX = CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A = CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B = CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D = CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_BMUX = CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_CMUX = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A = CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_AMUX = CLBLM_R_X5Y124_SLICE_X7Y124_A5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_BMUX = CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_DMUX = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A = CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B = CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_AMUX = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CMUX = CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A = CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_AMUX = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_AMUX = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_DMUX = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A = CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B = CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_DMUX = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A = CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B = CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A = CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B = CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_AMUX = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CMUX = CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A = CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B = CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C = CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A = CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_AMUX = CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_BMUX = CLBLM_R_X5Y129_SLICE_X6Y129_BO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A = CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B = CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_AMUX = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_BMUX = CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_CMUX = CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_CMUX = CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_AMUX = CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B = CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_DMUX = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CMUX = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_AMUX = CLBLM_R_X7Y119_SLICE_X9Y119_A5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_BMUX = CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CMUX = CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_DMUX = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CMUX = CLBLM_R_X7Y121_SLICE_X9Y121_C5Q;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_DMUX = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_BMUX = CLBLM_R_X7Y122_SLICE_X8Y122_B5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A = CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_BMUX = CLBLM_R_X7Y122_SLICE_X9Y122_B5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A = CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B = CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C = CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CMUX = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_DMUX = CLBLM_R_X7Y123_SLICE_X8Y123_DO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A = CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B = CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_DMUX = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A = CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B = CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A = CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C = CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_DMUX = CLBLM_R_X7Y125_SLICE_X9Y125_D5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_AMUX = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A = CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D = CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_CMUX = CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A = CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B = CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C = CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D = CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A = CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C = CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_AMUX = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D = CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_AMUX = CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_CMUX = CLBLM_R_X11Y115_SLICE_X15Y115_CO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A = CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_AMUX = CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_BMUX = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A = CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A = CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B = CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C = CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_AMUX = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_BMUX = CLBLM_R_X11Y118_SLICE_X14Y118_B5Q;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A = CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_AMUX = CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_BMUX = CLBLM_R_X11Y119_SLICE_X15Y119_B5Q;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_DMUX = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_CMUX = CLBLM_R_X11Y120_SLICE_X14Y120_CO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A = CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B = CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C = CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_BMUX = CLBLM_R_X11Y120_SLICE_X15Y120_B5Q;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_AMUX = CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_BMUX = CLBLM_R_X11Y121_SLICE_X14Y121_B5Q;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A = CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_AMUX = CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_BMUX = CLBLM_R_X11Y122_SLICE_X14Y122_BO5;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B = CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_DMUX = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A = CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B = CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C = CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_CMUX = CLBLM_R_X11Y124_SLICE_X14Y124_C5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_DMUX = CLBLM_R_X11Y124_SLICE_X14Y124_D5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A = CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_AMUX = CLBLM_R_X11Y124_SLICE_X15Y124_A5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_CMUX = CLBLM_R_X11Y124_SLICE_X15Y124_C5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A = CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C = CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A = CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B = CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C = CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C = CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D = CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_AMUX = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_BMUX = CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A = CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B = CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_BMUX = CLBLM_R_X11Y126_SLICE_X15Y126_BO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_CMUX = CLBLM_R_X11Y126_SLICE_X15Y126_CO5;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A = CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D = CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_CMUX = CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A = CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A = CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B = CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A = CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B = CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C = CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A = CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B = CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C = CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D = CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A = CLBLM_R_X13Y116_SLICE_X18Y116_AO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B = CLBLM_R_X13Y116_SLICE_X18Y116_BO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C = CLBLM_R_X13Y116_SLICE_X18Y116_CO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D = CLBLM_R_X13Y116_SLICE_X18Y116_DO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_BMUX = CLBLM_R_X13Y116_SLICE_X18Y116_BO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A = CLBLM_R_X13Y116_SLICE_X19Y116_AO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B = CLBLM_R_X13Y116_SLICE_X19Y116_BO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C = CLBLM_R_X13Y116_SLICE_X19Y116_CO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D = CLBLM_R_X13Y116_SLICE_X19Y116_DO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A = CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B = CLBLM_R_X13Y117_SLICE_X18Y117_BO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C = CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D = CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_AMUX = CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A = CLBLM_R_X13Y117_SLICE_X19Y117_AO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B = CLBLM_R_X13Y117_SLICE_X19Y117_BO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C = CLBLM_R_X13Y117_SLICE_X19Y117_CO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D = CLBLM_R_X13Y117_SLICE_X19Y117_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A = CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B = CLBLM_R_X13Y118_SLICE_X18Y118_BO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C = CLBLM_R_X13Y118_SLICE_X18Y118_CO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D = CLBLM_R_X13Y118_SLICE_X18Y118_DO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A = CLBLM_R_X13Y118_SLICE_X19Y118_AO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B = CLBLM_R_X13Y118_SLICE_X19Y118_BO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C = CLBLM_R_X13Y118_SLICE_X19Y118_CO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D = CLBLM_R_X13Y118_SLICE_X19Y118_DO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A = CLBLM_R_X13Y119_SLICE_X18Y119_AO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B = CLBLM_R_X13Y119_SLICE_X18Y119_BO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C = CLBLM_R_X13Y119_SLICE_X18Y119_CO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D = CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_AMUX = CLBLM_R_X13Y119_SLICE_X18Y119_A5Q;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_BMUX = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A = CLBLM_R_X13Y119_SLICE_X19Y119_AO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B = CLBLM_R_X13Y119_SLICE_X19Y119_BO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C = CLBLM_R_X13Y119_SLICE_X19Y119_CO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D = CLBLM_R_X13Y119_SLICE_X19Y119_DO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A = CLBLM_R_X13Y120_SLICE_X18Y120_AO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B = CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_CMUX = CLBLM_R_X13Y120_SLICE_X18Y120_CO5;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_DMUX = CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A = CLBLM_R_X13Y120_SLICE_X19Y120_AO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B = CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C = CLBLM_R_X13Y120_SLICE_X19Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D = CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_AMUX = CLBLM_R_X13Y120_SLICE_X19Y120_A5Q;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_BMUX = CLBLM_R_X13Y120_SLICE_X19Y120_BO5;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A = CLBLM_R_X13Y121_SLICE_X18Y121_AO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B = CLBLM_R_X13Y121_SLICE_X18Y121_BO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C = CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A = CLBLM_R_X13Y121_SLICE_X19Y121_AO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B = CLBLM_R_X13Y121_SLICE_X19Y121_BO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C = CLBLM_R_X13Y121_SLICE_X19Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D = CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A = CLBLM_R_X13Y122_SLICE_X18Y122_AO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B = CLBLM_R_X13Y122_SLICE_X18Y122_BO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D = CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A = CLBLM_R_X13Y122_SLICE_X19Y122_AO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B = CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C = CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D = CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A = CLBLM_R_X13Y123_SLICE_X18Y123_AO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B = CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C = CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D = CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A = CLBLM_R_X13Y123_SLICE_X19Y123_AO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B = CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C = CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D = CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A = CLBLM_R_X13Y124_SLICE_X18Y124_AO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B = CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C = CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D = CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A = CLBLM_R_X13Y124_SLICE_X19Y124_AO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B = CLBLM_R_X13Y124_SLICE_X19Y124_BO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C = CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D = CLBLM_R_X13Y124_SLICE_X19Y124_DO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_CMUX = CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A = CLBLM_R_X13Y125_SLICE_X18Y125_AO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C = CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D = CLBLM_R_X13Y125_SLICE_X18Y125_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_BMUX = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_CMUX = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_DMUX = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A = CLBLM_R_X13Y125_SLICE_X19Y125_AO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C = CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D = CLBLM_R_X13Y125_SLICE_X19Y125_DO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_BMUX = CLBLM_R_X13Y125_SLICE_X19Y125_BO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B = CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C = CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_AMUX = CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_BMUX = CLBLM_R_X13Y126_SLICE_X18Y126_BO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_DMUX = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A = CLBLM_R_X13Y126_SLICE_X19Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B = CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C = CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D = CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D = CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A = CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B = CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C = CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B = CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D = CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_A = CLBLM_R_X25Y143_SLICE_X36Y143_AO6;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_B = CLBLM_R_X25Y143_SLICE_X36Y143_BO6;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_C = CLBLM_R_X25Y143_SLICE_X36Y143_CO6;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_D = CLBLM_R_X25Y143_SLICE_X36Y143_DO6;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_AMUX = CLBLM_R_X25Y143_SLICE_X36Y143_AO5;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_A = CLBLM_R_X25Y143_SLICE_X37Y143_AO6;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_B = CLBLM_R_X25Y143_SLICE_X37Y143_BO6;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_C = CLBLM_R_X25Y143_SLICE_X37Y143_CO6;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_D = CLBLM_R_X25Y143_SLICE_X37Y143_DO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B = CLBLM_R_X37Y120_SLICE_X56Y120_BO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C = CLBLM_R_X37Y120_SLICE_X56Y120_CO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D = CLBLM_R_X37Y120_SLICE_X56Y120_DO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A = CLBLM_R_X37Y120_SLICE_X57Y120_AO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B = CLBLM_R_X37Y120_SLICE_X57Y120_BO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C = CLBLM_R_X37Y120_SLICE_X57Y120_CO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D = CLBLM_R_X37Y120_SLICE_X57Y120_DO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A = CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B = CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C = CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D = CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B = CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C = CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D = CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_AMUX = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A = CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B = CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C = CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D = CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B = CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C = CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D = CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_AMUX = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A = CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B = CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C = CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D = CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B = CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C = CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D = CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_AMUX = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_L_X12Y117_SLICE_X16Y117_D5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_L_X12Y117_SLICE_X16Y117_DQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_R_X5Y122_SLICE_X6Y122_B5Q;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X8Y126_SLICE_X11Y126_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X7Y122_SLICE_X8Y122_B5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X7Y121_SLICE_X9Y121_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y118_SLICE_X3Y118_A5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X13Y118_SLICE_X19Y118_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X25Y143_SLICE_X36Y143_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X25Y143_SLICE_X36Y143_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D4 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B6 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_AX = CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = CLBLM_R_X3Y120_SLICE_X3Y120_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = CLBLM_R_X3Y120_SLICE_X3Y120_A5Q;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = CLBLL_L_X4Y119_SLICE_X5Y119_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A1 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A2 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A4 = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A5 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B1 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B3 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B4 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_BX = CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D6 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B5 = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C4 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D4 = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D6 = 1'b1;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_A5 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_AX = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = CLBLM_R_X3Y120_SLICE_X3Y120_A5Q;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_AX = CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C3 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C1 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A3 = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A4 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C6 = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D6 = 1'b1;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A1 = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A5 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_A5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_A6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B1 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B2 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B3 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B4 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B5 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D2 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D3 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C1 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C3 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C4 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C5 = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C6 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D5 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D2 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D4 = CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D6 = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_B3 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_B4 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_B5 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_B6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B5 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B6 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_C4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C3 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_C5 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C5 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A2 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A3 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A5 = CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A6 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_D4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C6 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_D5 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_D6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D6 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A3 = CLBLM_L_X12Y116_SLICE_X16Y116_AO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A4 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A5 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A6 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B1 = CLBLM_L_X12Y116_SLICE_X16Y116_AO5;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B2 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B4 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B5 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C3 = CLBLM_R_X13Y117_SLICE_X19Y117_BQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C4 = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A2 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A6 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D1 = CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D2 = CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D3 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D4 = CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D5 = CLBLM_R_X13Y116_SLICE_X18Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D6 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C2 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A1 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A2 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A3 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A4 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A5 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C5 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_AX = CLBLM_L_X12Y117_SLICE_X16Y117_DQ;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C6 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B3 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B4 = CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B5 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B6 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D3 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C2 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C3 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C4 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C5 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C6 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A2 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A6 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D2 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D3 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D4 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D5 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B3 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_SR = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A6 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A1 = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A2 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A3 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A4 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A5 = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B1 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B2 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B3 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B4 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B5 = CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B6 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C1 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C2 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C3 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C4 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C5 = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D1 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D3 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D4 = CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D5 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A1 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A3 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A4 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A5 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A6 = CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C6 = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A1 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A3 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A4 = CLBLM_R_X11Y118_SLICE_X14Y118_B5Q;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B1 = CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B2 = CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B3 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B4 = CLBLM_L_X12Y117_SLICE_X16Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B5 = CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C2 = CLBLM_R_X13Y117_SLICE_X18Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C3 = CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C4 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C5 = CLBLM_L_X12Y117_SLICE_X17Y117_BO5;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C6 = CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D1 = CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D2 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D4 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D5 = CLBLM_R_X13Y116_SLICE_X18Y116_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D6 = CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A2 = CLBLM_L_X12Y117_SLICE_X16Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A3 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A4 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A5 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A6 = CLBLM_L_X12Y118_SLICE_X16Y118_CQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B1 = CLBLM_R_X13Y118_SLICE_X18Y118_DQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B2 = CLBLM_L_X12Y117_SLICE_X16Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B6 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C2 = CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C4 = CLBLM_L_X12Y117_SLICE_X16Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C5 = CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D3 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D4 = CLBLM_R_X13Y118_SLICE_X18Y118_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D5 = CLBLM_R_X11Y118_SLICE_X14Y118_B5Q;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A2 = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B6 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A5 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B3 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B5 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B6 = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C1 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C2 = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C3 = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C4 = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C5 = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C6 = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D2 = CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D3 = CLBLM_L_X10Y123_SLICE_X12Y123_C5Q;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D5 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A1 = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A2 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A3 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A4 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A5 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A6 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B1 = CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B5 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B6 = CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C1 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C2 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C3 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C4 = CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C6 = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A1 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A3 = CLBLM_L_X12Y118_SLICE_X17Y118_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A4 = CLBLM_R_X13Y118_SLICE_X18Y118_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B5 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B6 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C1 = CLBLM_R_X13Y118_SLICE_X18Y118_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C2 = CLBLM_R_X13Y117_SLICE_X19Y117_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C3 = CLBLM_R_X13Y118_SLICE_X18Y118_DQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C5 = CLBLM_L_X12Y118_SLICE_X17Y118_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C6 = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D1 = CLBLM_R_X11Y118_SLICE_X14Y118_CQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D2 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D3 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A1 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A2 = CLBLM_L_X12Y118_SLICE_X16Y118_DQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A3 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A5 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B1 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B2 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B5 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B6 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C2 = CLBLM_L_X12Y118_SLICE_X16Y118_CQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C3 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C4 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C6 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D2 = CLBLM_L_X12Y119_SLICE_X17Y119_BQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D3 = CLBLM_L_X12Y118_SLICE_X16Y118_DQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D4 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B4 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B6 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C5 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C6 = CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C2 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B2 = CLBLM_R_X25Y143_SLICE_X36Y143_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B3 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B4 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B5 = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B6 = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D5 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C1 = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C3 = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C4 = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C5 = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C6 = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A1 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C4 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D1 = CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D2 = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D3 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D4 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D5 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D6 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_AX = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A1 = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A3 = CLBLM_L_X12Y119_SLICE_X17Y119_AQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A5 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B5 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_AX = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_D5Q;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B1 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B2 = CLBLM_L_X12Y119_SLICE_X17Y119_BQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B5 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B6 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = CLBLL_L_X4Y120_SLICE_X4Y120_DQ;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C2 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C4 = CLBLM_L_X12Y119_SLICE_X17Y119_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C5 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C6 = CLBLM_L_X12Y118_SLICE_X17Y118_BQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = CLBLL_L_X4Y120_SLICE_X4Y120_A5Q;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D1 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D2 = CLBLM_L_X12Y119_SLICE_X17Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D3 = CLBLM_R_X13Y121_SLICE_X18Y121_DQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D4 = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D5 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D6 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A1 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_BX = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A3 = CLBLM_L_X12Y119_SLICE_X16Y119_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A4 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A5 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A6 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B2 = CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B4 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B6 = CLBLL_L_X4Y120_SLICE_X4Y120_DQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C4 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C1 = CLBLM_R_X13Y120_SLICE_X19Y120_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C2 = CLBLM_L_X12Y119_SLICE_X16Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C3 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = CLBLL_L_X4Y119_SLICE_X5Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C6 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D2 = CLBLM_L_X12Y119_SLICE_X16Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D3 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D6 = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A1 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B2 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = CLBLL_L_X4Y120_SLICE_X4Y120_DQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = CLBLM_L_X12Y116_SLICE_X17Y116_CQ;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B2 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D5 = CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D6 = CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D6 = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A1 = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A2 = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A3 = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A4 = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A5 = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A6 = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B1 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B2 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B3 = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B4 = CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B5 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B6 = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C1 = CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C2 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C3 = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C4 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D1 = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D2 = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D3 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D4 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D6 = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A1 = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A2 = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A3 = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A4 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A5 = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A6 = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B2 = CLBLM_R_X25Y143_SLICE_X36Y143_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B4 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C1 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C2 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C3 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C4 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C5 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D1 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D2 = CLBLM_R_X25Y143_SLICE_X36Y143_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D3 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D4 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D5 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D6 = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A2 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A3 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A4 = CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A6 = CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B1 = CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B3 = CLBLM_L_X10Y120_SLICE_X12Y120_A5Q;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C1 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C2 = CLBLM_L_X12Y120_SLICE_X17Y120_CQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C3 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D1 = CLBLM_L_X12Y119_SLICE_X17Y119_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D2 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D3 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D4 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D5 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A3 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A5 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A6 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B2 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B3 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B4 = CLBLM_R_X13Y118_SLICE_X18Y118_DQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B6 = CLBLM_L_X10Y123_SLICE_X12Y123_DQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C1 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C2 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C3 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C4 = CLBLM_L_X12Y120_SLICE_X17Y120_CQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C6 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D1 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D2 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D3 = CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D6 = CLBLM_L_X10Y123_SLICE_X12Y123_DQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C2 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B5 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C1 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C2 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D3 = CLBLM_R_X3Y127_SLICE_X3Y127_AO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D4 = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D5 = CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A6 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B1 = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B2 = CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B3 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B5 = CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B6 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C3 = CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C6 = CLBLM_R_X25Y143_SLICE_X36Y143_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A1 = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A3 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A5 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B2 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B4 = CLBLM_L_X12Y121_SLICE_X17Y121_DO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B5 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B6 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C3 = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C5 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C6 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D1 = CLBLM_L_X12Y119_SLICE_X17Y119_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D2 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D3 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D4 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D5 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A2 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A3 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A4 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A5 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_AX = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B1 = CLBLM_L_X12Y123_SLICE_X16Y123_DQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B2 = CLBLM_L_X12Y116_SLICE_X17Y116_CQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B3 = CLBLM_L_X12Y120_SLICE_X17Y120_CQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D1 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C1 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C2 = CLBLM_L_X12Y121_SLICE_X16Y121_CQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C4 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D4 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D5 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A2 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A4 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B1 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B2 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B3 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B4 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C1 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C2 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C3 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C4 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D1 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D2 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D3 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D4 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B1 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B2 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B3 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B4 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C1 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C2 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C3 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C4 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D1 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D2 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D3 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D4 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A1 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A2 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A3 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A4 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A5 = CLBLM_R_X11Y122_SLICE_X15Y122_DQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_AX = CLBLM_R_X11Y122_SLICE_X15Y122_DQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B1 = CLBLM_L_X12Y122_SLICE_X16Y122_DQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B2 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B4 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B5 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C1 = CLBLM_L_X12Y121_SLICE_X16Y121_CQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C2 = CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C3 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C4 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C5 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D1 = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D2 = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D3 = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D4 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D5 = CLBLM_R_X11Y122_SLICE_X15Y122_CQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D6 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_SR = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A1 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A2 = CLBLM_L_X12Y122_SLICE_X16Y122_DQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A5 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B2 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B4 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B6 = CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C2 = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C3 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C4 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C5 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C6 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D2 = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D4 = CLBLM_L_X12Y122_SLICE_X16Y122_DQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D5 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A2 = CLBLM_R_X11Y120_SLICE_X14Y120_DQ;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A4 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A5 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A1 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A2 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A4 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B2 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B4 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B2 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C1 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C2 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C4 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B4 = CLBLM_L_X8Y115_SLICE_X11Y115_DQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D1 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D2 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D4 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A1 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A3 = CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A4 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B1 = CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B2 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B3 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B4 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B5 = CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B6 = CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C1 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C2 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C4 = CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C6 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C4 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D1 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D2 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D4 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D1 = CLBLL_L_X4Y121_SLICE_X5Y121_DQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D2 = CLBLM_L_X8Y115_SLICE_X11Y115_CQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A1 = CLBLM_L_X10Y125_SLICE_X13Y125_DQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A2 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A3 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B1 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B3 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B4 = CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B5 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B6 = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A6 = CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C2 = CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C3 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B1 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B2 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D1 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C3 = CLBLM_L_X8Y116_SLICE_X11Y116_C5Q;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C5 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D3 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D4 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A1 = CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A3 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A4 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A5 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D6 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A6 = CLBLM_R_X13Y122_SLICE_X18Y122_CQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B1 = CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B2 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B3 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A1 = CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A3 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A4 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A5 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C2 = CLBLM_L_X12Y123_SLICE_X16Y123_CQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B3 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B4 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D1 = CLBLM_R_X13Y119_SLICE_X19Y119_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C6 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D6 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B4 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A3 = CLBLM_R_X13Y117_SLICE_X19Y117_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A4 = CLBLM_R_X13Y117_SLICE_X19Y117_CQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A5 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B2 = CLBLM_R_X13Y117_SLICE_X19Y117_BQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B3 = CLBLM_R_X13Y117_SLICE_X19Y117_AQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B4 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C1 = CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C2 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C6 = CLBLM_R_X13Y117_SLICE_X19Y117_CQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A1 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A2 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A3 = CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A5 = CLBLM_R_X13Y117_SLICE_X19Y117_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A6 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B1 = CLBLM_R_X13Y118_SLICE_X18Y118_CQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B3 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B4 = CLBLM_R_X13Y118_SLICE_X18Y118_DQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B5 = CLBLM_R_X13Y117_SLICE_X19Y117_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B6 = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C1 = CLBLM_R_X13Y119_SLICE_X19Y119_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C2 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C3 = CLBLM_L_X12Y117_SLICE_X16Y117_BQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C5 = CLBLM_R_X13Y118_SLICE_X18Y118_CQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D1 = CLBLM_R_X13Y119_SLICE_X19Y119_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D2 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D3 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D6 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A1 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A2 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A3 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A5 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A6 = CLBLM_L_X12Y118_SLICE_X17Y118_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B3 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B4 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B1 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B2 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B3 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B5 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B6 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A1 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A2 = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A3 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A4 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A5 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A6 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C1 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C2 = CLBLM_L_X12Y123_SLICE_X17Y123_CQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B2 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B4 = CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B5 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B6 = CLBLM_L_X8Y116_SLICE_X11Y116_C5Q;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D1 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D2 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C1 = CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C2 = CLBLM_L_X12Y115_SLICE_X16Y115_BO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C3 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C4 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C5 = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D3 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D4 = CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D5 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D6 = CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A2 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A3 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D1 = CLBLM_R_X11Y115_SLICE_X15Y115_CO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D2 = CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D3 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D4 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D5 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C3 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C5 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A1 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A3 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A4 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A6 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C6 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B2 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B3 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B4 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B5 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C1 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C3 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C4 = CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D2 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D4 = CLBLM_L_X8Y116_SLICE_X11Y116_C5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D5 = CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A3 = CLBLM_R_X13Y118_SLICE_X19Y118_AQ;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A6 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A2 = CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A3 = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A5 = CLBLM_R_X13Y118_SLICE_X19Y118_AQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B2 = CLBLM_R_X13Y118_SLICE_X18Y118_BQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B3 = CLBLM_R_X13Y122_SLICE_X18Y122_CQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B4 = CLBLM_R_X13Y117_SLICE_X19Y117_BQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C1 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C2 = CLBLM_R_X13Y118_SLICE_X18Y118_CQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C4 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D2 = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D3 = CLBLM_R_X13Y118_SLICE_X18Y118_DQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D5 = CLBLM_L_X10Y118_SLICE_X12Y118_DQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A3 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A4 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A1 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A2 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A3 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A4 = CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A6 = CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A5 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B1 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B2 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B3 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B4 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B5 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B6 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_DQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C2 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C3 = CLBLM_L_X10Y125_SLICE_X13Y125_DQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C4 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C5 = CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C6 = CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A2 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A3 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A4 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A5 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B2 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D1 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D2 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B4 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B5 = CLBLM_L_X8Y115_SLICE_X11Y115_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B6 = CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C1 = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C2 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C3 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C4 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C6 = CLBLM_R_X11Y124_SLICE_X14Y124_D5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A1 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A2 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A3 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A5 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A6 = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D1 = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D2 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D3 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D4 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D5 = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B3 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B5 = CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D6 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B1 = CLBLM_L_X12Y126_SLICE_X16Y126_AO5;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B2 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A1 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C2 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C3 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C5 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C6 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A2 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A3 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A4 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A5 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A6 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C1 = CLBLM_L_X8Y117_SLICE_X11Y117_CO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C3 = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C4 = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C5 = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C6 = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D3 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D6 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D6 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A1 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A3 = CLBLM_R_X13Y119_SLICE_X19Y119_AQ;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A6 = CLBLM_R_X13Y118_SLICE_X18Y118_CQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B3 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B4 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B5 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B6 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C2 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C3 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C4 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C5 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C6 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D2 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D3 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D4 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D5 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D6 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A1 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A2 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A3 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A4 = CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A5 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_AX = CLBLM_R_X13Y119_SLICE_X18Y119_BO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B1 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B2 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B3 = CLBLM_L_X8Y117_SLICE_X10Y117_A5Q;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B5 = CLBLM_R_X13Y119_SLICE_X18Y119_A5Q;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C1 = CLBLM_L_X12Y118_SLICE_X17Y118_BQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C2 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C3 = CLBLM_L_X10Y123_SLICE_X13Y123_C5Q;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C4 = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D1 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D2 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D3 = CLBLM_L_X12Y123_SLICE_X16Y123_DQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D4 = CLBLM_L_X12Y118_SLICE_X17Y118_BQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D5 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D6 = CLBLM_R_X13Y119_SLICE_X19Y119_BQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A1 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A2 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A3 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B2 = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B3 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B4 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B5 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B6 = CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C1 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C2 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C3 = CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C4 = CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A2 = CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A3 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A4 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A6 = CLBLM_L_X8Y115_SLICE_X11Y115_CQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B1 = CLBLM_R_X11Y124_SLICE_X14Y124_DQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B2 = CLBLM_L_X12Y119_SLICE_X17Y119_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B3 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B4 = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B5 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B6 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C1 = CLBLM_L_X12Y119_SLICE_X17Y119_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C2 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C3 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_C5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C5 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C6 = CLBLM_L_X12Y118_SLICE_X16Y118_DQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D5 = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A1 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A2 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A3 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A4 = CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A5 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D3 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D4 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D5 = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D6 = CLBLM_L_X12Y119_SLICE_X17Y119_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B4 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B5 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B1 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_BX = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B2 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C1 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C2 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C3 = CLBLM_R_X11Y126_SLICE_X15Y126_BO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C4 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C5 = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C6 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A2 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A4 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A5 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B1 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D2 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D4 = CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B3 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B5 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C2 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C4 = CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C5 = CLBLM_R_X13Y119_SLICE_X19Y119_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_SR = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D1 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D3 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D5 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A2 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A3 = CLBLM_R_X13Y120_SLICE_X19Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A4 = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_AX = CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B2 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B3 = CLBLM_R_X13Y120_SLICE_X19Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B4 = CLBLM_R_X13Y118_SLICE_X18Y118_CQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B6 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C1 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C2 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C3 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C4 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C5 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C6 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D1 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D2 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D3 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D4 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D5 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D6 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A1 = CLBLM_R_X13Y121_SLICE_X18Y121_CQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A3 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A4 = CLBLM_R_X13Y117_SLICE_X19Y117_CQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A5 = CLBLM_R_X13Y120_SLICE_X18Y120_CO5;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A6 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B1 = CLBLM_R_X13Y120_SLICE_X19Y120_A5Q;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B2 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B4 = CLBLM_L_X12Y120_SLICE_X17Y120_BO5;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B5 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C1 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C2 = CLBLM_R_X13Y119_SLICE_X18Y119_A5Q;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C4 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C5 = CLBLM_R_X13Y120_SLICE_X19Y120_A5Q;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C6 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D1 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D2 = CLBLM_R_X13Y119_SLICE_X18Y119_A5Q;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D3 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D4 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D5 = CLBLM_R_X13Y121_SLICE_X18Y121_CQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A2 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A3 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B2 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B3 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C2 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A6 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A3 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D2 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D3 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C1 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C2 = CLBLM_L_X8Y117_SLICE_X10Y117_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A1 = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A2 = CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A3 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A4 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B2 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B3 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D5 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D6 = CLBLM_R_X11Y124_SLICE_X14Y124_D5Q;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C2 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C3 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A5 = CLBLM_R_X13Y119_SLICE_X19Y119_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A6 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B1 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C1 = CLBLM_L_X8Y117_SLICE_X11Y117_CO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C5 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C6 = CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C2 = CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C3 = CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D4 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D5 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D1 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A1 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A6 = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A1 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A3 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A4 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A5 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B1 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B3 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B4 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B5 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D3 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C3 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C4 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B3 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D1 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D3 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D4 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D5 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A1 = CLBLM_R_X13Y121_SLICE_X18Y121_CQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A3 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A4 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A6 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B2 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B5 = CLBLM_L_X12Y118_SLICE_X17Y118_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B6 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C1 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C2 = CLBLM_R_X13Y121_SLICE_X18Y121_CQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C3 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C4 = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C6 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C3 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C4 = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D1 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D3 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D6 = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D4 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C6 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_L_X12Y117_SLICE_X16Y117_D5Q;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A1 = CLBLM_L_X12Y123_SLICE_X16Y123_DQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A2 = CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A4 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A5 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B1 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B3 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B4 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B5 = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C1 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C2 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C3 = CLBLM_R_X11Y124_SLICE_X14Y124_DQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C5 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D1 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D2 = CLBLM_L_X8Y118_SLICE_X11Y118_CQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D3 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D4 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A3 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A4 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A6 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B3 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B4 = CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B5 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B6 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_AX = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C2 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D3 = CLBLM_L_X10Y118_SLICE_X12Y118_DQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D5 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D6 = CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D5 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A2 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A3 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A4 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B1 = CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B2 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B3 = CLBLM_R_X11Y122_SLICE_X15Y122_DQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B4 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B5 = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B6 = CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C1 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C2 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C3 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C4 = CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C5 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C6 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D1 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D2 = CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D3 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D4 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D5 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D6 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A1 = CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A2 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A4 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A5 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A6 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B1 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B2 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B4 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B5 = CLBLM_R_X13Y119_SLICE_X19Y119_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B6 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C1 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C2 = CLBLM_R_X13Y122_SLICE_X18Y122_CQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C4 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C6 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D1 = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D2 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D3 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D4 = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D5 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D6 = 1'b1;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C6 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B5 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A2 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A3 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A4 = CLBLM_L_X12Y118_SLICE_X16Y118_DQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A6 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C1 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B1 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B2 = CLBLM_L_X12Y119_SLICE_X17Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B3 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B4 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B5 = CLBLM_L_X12Y118_SLICE_X16Y118_DQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B6 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C2 = CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C3 = CLBLM_R_X5Y122_SLICE_X6Y122_A5Q;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C1 = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C2 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C3 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C4 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C5 = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C6 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C6 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D2 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D4 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D6 = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A1 = CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A3 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A4 = CLBLM_R_X13Y119_SLICE_X18Y119_A5Q;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A6 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A3 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B2 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B4 = CLBLM_L_X10Y116_SLICE_X12Y116_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A4 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C1 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C2 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C5 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C6 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A6 = 1'b1;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D3 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D5 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D6 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_A1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_A2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_A3 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_A4 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_A6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B1 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_B1 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_B2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_B3 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_B4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_B5 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_B6 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_C1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B3 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_C2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_C3 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_C4 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_C5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B4 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_C6 = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_D1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B5 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_D2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_D3 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_D4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A2 = CLBLM_L_X12Y123_SLICE_X17Y123_CQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A3 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_D5 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B1 = CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B2 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B4 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B5 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B6 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_A3 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_A4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C1 = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C2 = CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C3 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C4 = CLBLM_L_X12Y123_SLICE_X16Y123_DQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C6 = CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_B1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_B2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_C1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C1 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_C2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_C3 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D1 = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C2 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D2 = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D3 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D4 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D5 = CLBLM_R_X13Y124_SLICE_X19Y124_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C3 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D6 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_C6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C4 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_D1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A1 = CLBLM_R_X13Y125_SLICE_X18Y125_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A2 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A3 = CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C5 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A4 = CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A6 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_D2 = 1'b1;
  assign CLBLM_R_X25Y143_SLICE_X36Y143_D3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B1 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B2 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B3 = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B2 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B5 = CLBLM_R_X13Y124_SLICE_X18Y124_AO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X7Y122_SLICE_X8Y122_B5Q;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C1 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C2 = CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C3 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C4 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C5 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C6 = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D2 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D3 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D5 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D2 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D3 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D5 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C4 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B4 = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C5 = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C6 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_C5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A1 = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A3 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A6 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B1 = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B2 = CLBLM_L_X10Y119_SLICE_X12Y119_B5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B3 = CLBLM_L_X10Y120_SLICE_X12Y120_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B4 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B5 = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B6 = CLBLM_R_X7Y122_SLICE_X9Y122_B5Q;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C1 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C2 = CLBLM_L_X10Y123_SLICE_X13Y123_C5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C3 = CLBLM_L_X12Y123_SLICE_X16Y123_DQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C5 = CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C6 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D2 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A3 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_DQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D3 = CLBLM_R_X11Y120_SLICE_X15Y120_DQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D4 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B3 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B5 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D5 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D5 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A2 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A3 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A5 = CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B4 = CLBLM_L_X10Y119_SLICE_X12Y119_B5Q;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B6 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_BX = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C1 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C5 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B2 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A4 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D1 = CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D2 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D5 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D6 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B3 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B5 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A1 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A2 = CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A3 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A4 = CLBLM_L_X12Y123_SLICE_X17Y123_CQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A5 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A6 = CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B2 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B3 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B4 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B5 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B6 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C1 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C2 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C3 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B5 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C5 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B6 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A1 = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A2 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A3 = CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A4 = CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B1 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B2 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B3 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A1 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A2 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A4 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A5 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C1 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C2 = CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D1 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D2 = CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D3 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C2 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C6 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C5 = CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D4 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D6 = CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C4 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_AX = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A1 = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A3 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A6 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B1 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B2 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B3 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B4 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B5 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B2 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C1 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C2 = CLBLL_L_X4Y120_SLICE_X5Y120_DQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C3 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C4 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C6 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D2 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D4 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A2 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A4 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A6 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B1 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_C5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = CLBLM_R_X3Y118_SLICE_X3Y118_A5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B5 = CLBLM_L_X12Y123_SLICE_X16Y123_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B6 = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C1 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C2 = CLBLM_L_X12Y123_SLICE_X16Y123_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C3 = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C4 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C5 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D1 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_B5Q;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D4 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D5 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D6 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A1 = CLBLM_R_X13Y125_SLICE_X19Y125_DO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A2 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A5 = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A6 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_C5Q;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B2 = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B3 = CLBLM_R_X13Y124_SLICE_X19Y124_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A2 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A3 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A4 = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A5 = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A6 = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C1 = CLBLM_R_X13Y122_SLICE_X18Y122_CQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C2 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B1 = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B2 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B3 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B4 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D5 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C1 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C2 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C3 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D6 = CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A2 = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A3 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D1 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D2 = CLBLM_R_X11Y124_SLICE_X14Y124_D5Q;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D3 = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D4 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_C5Q;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B1 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B2 = CLBLM_R_X13Y125_SLICE_X19Y125_BO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B3 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A1 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A2 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A3 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A4 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A5 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C1 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B1 = CLBLM_R_X11Y121_SLICE_X14Y121_B5Q;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B6 = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D1 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C1 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C2 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C3 = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C4 = CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C5 = CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C6 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D2 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D3 = CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D2 = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D3 = CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D5 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D6 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A2 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A3 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A4 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A5 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_AX = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B2 = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B3 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B5 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B6 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C1 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C4 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C6 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A2 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A3 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A4 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A5 = CLBLM_L_X12Y117_SLICE_X16Y117_D5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D1 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D4 = CLBLM_R_X11Y121_SLICE_X15Y121_DQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B2 = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B4 = CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C1 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C2 = CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A1 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A2 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A3 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A6 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C3 = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C4 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B2 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B3 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B4 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B5 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_C5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D3 = CLBLM_R_X3Y118_SLICE_X3Y118_A5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D4 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D5 = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C1 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C3 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D2 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D4 = CLBLM_R_X7Y122_SLICE_X9Y122_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A5 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A6 = CLBLL_L_X4Y119_SLICE_X5Y119_A5Q;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B1 = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B2 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B4 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B5 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B6 = CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C1 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C3 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C4 = CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C5 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C6 = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A3 = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A2 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A3 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A4 = CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D1 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D2 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D4 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A5 = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A6 = CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A1 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A2 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A4 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A5 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B3 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B4 = CLBLM_L_X8Y123_SLICE_X11Y123_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B2 = CLBLM_L_X10Y120_SLICE_X12Y120_A5Q;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B6 = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C1 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C2 = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C3 = CLBLM_R_X11Y116_SLICE_X15Y116_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C4 = CLBLM_L_X12Y119_SLICE_X17Y119_A5Q;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C5 = CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C6 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A1 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A2 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A3 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D1 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D2 = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D3 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D4 = CLBLM_L_X12Y116_SLICE_X17Y116_CQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D5 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D6 = CLBLM_R_X11Y124_SLICE_X14Y124_DQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A5 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B1 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B2 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B3 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A1 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A3 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A5 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A6 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C1 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C2 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B1 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B2 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C1 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B3 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B6 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C2 = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D1 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C3 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C5 = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C4 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C6 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D4 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D6 = CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D4 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D2 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D3 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D4 = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D5 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A1 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A2 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A3 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A6 = CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B2 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B4 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B5 = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C1 = CLBLM_L_X10Y123_SLICE_X13Y123_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C3 = CLBLM_L_X10Y123_SLICE_X13Y123_DQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C4 = CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D2 = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = CLBLL_L_X4Y120_SLICE_X4Y120_CQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A1 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A3 = CLBLM_L_X10Y124_SLICE_X12Y124_C5Q;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A4 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B3 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B5 = CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B6 = CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C4 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C5 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C2 = CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D1 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = CLBLM_R_X5Y118_SLICE_X6Y118_DQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D6 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_AX = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = CLBLM_L_X8Y116_SLICE_X11Y116_CQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B4 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = CLBLL_L_X4Y119_SLICE_X5Y119_DQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B6 = CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = CLBLL_L_X4Y119_SLICE_X5Y119_DQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B1 = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A2 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A4 = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A6 = CLBLM_L_X12Y118_SLICE_X16Y118_CQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C2 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B1 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B4 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B5 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B6 = CLBLM_L_X12Y118_SLICE_X16Y118_CQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D2 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C1 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C2 = CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C3 = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C4 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D4 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A2 = CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A3 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A5 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A6 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D1 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D2 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D3 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D4 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D6 = CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A1 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A2 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A3 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A4 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C3 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B4 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B5 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C1 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C2 = CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C4 = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D4 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D6 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D2 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D3 = CLBLM_R_X11Y117_SLICE_X14Y117_DQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B3 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B5 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B6 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A1 = CLBLM_L_X10Y125_SLICE_X13Y125_DQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A3 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A5 = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A6 = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C4 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B1 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B4 = CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B5 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C4 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C5 = CLBLM_R_X11Y120_SLICE_X15Y120_DQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A4 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A6 = CLBLM_L_X8Y116_SLICE_X11Y116_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D1 = CLBLM_R_X11Y124_SLICE_X15Y124_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D3 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D4 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = CLBLL_L_X4Y120_SLICE_X4Y120_CQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A2 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A6 = CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B2 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B3 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B4 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B5 = CLBLM_R_X11Y124_SLICE_X14Y124_D5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C2 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C4 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C5 = CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A1 = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D2 = CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D4 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D5 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D6 = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = CLBLL_L_X4Y121_SLICE_X5Y121_DQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = CLBLM_R_X11Y120_SLICE_X15Y120_B5Q;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = CLBLM_R_X5Y118_SLICE_X6Y118_DQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D2 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A2 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A3 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A6 = CLBLM_R_X11Y118_SLICE_X14Y118_CQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D3 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D4 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B1 = CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B2 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B3 = CLBLL_L_X4Y120_SLICE_X5Y120_DQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B4 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B5 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D5 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C1 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C2 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C3 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_AO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C5 = CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C6 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D2 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D3 = CLBLM_L_X12Y119_SLICE_X16Y119_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D4 = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D5 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D6 = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A1 = CLBLM_L_X10Y120_SLICE_X12Y120_B5Q;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A3 = CLBLM_L_X12Y119_SLICE_X16Y119_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A5 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B1 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B5 = CLBLM_R_X11Y119_SLICE_X15Y119_B5Q;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C5 = CLBLM_R_X13Y126_SLICE_X18Y126_BO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C3 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C2 = CLBLM_R_X11Y118_SLICE_X14Y118_CQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C4 = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C6 = CLBLL_L_X4Y121_SLICE_X5Y121_D5Q;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D1 = CLBLM_R_X13Y119_SLICE_X19Y119_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D3 = CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D4 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D5 = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D6 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C4 = 1'b1;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A1 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A2 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A3 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A5 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C5 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A6 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B4 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B5 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X8Y126_SLICE_X11Y126_A5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C3 = CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C4 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B1 = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C5 = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B2 = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C6 = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B3 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B4 = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A5 = CLBLM_L_X12Y125_SLICE_X16Y125_DQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A6 = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B5 = CLBLM_R_X7Y123_SLICE_X8Y123_DO5;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B6 = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C2 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A1 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B4 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B5 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B6 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A3 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A5 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C1 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C2 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C3 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C6 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B1 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B2 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D1 = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D2 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D3 = CLBLM_L_X12Y125_SLICE_X16Y125_DQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C2 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D6 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A1 = CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A2 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A4 = CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A5 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A6 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D1 = CLBLL_L_X4Y121_SLICE_X5Y121_D5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D2 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D5 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B4 = CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B5 = CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B6 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D6 = CLBLM_L_X8Y115_SLICE_X11Y115_DQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A2 = CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A3 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C4 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C5 = CLBLM_R_X11Y124_SLICE_X14Y124_C5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C6 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A6 = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B6 = CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D2 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D3 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D4 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D5 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C4 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C5 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C6 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_SR = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C1 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B2 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B3 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B6 = CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C1 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C3 = CLBLM_R_X7Y122_SLICE_X9Y122_B5Q;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D6 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C5 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C6 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D3 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D4 = CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D1 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D2 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D4 = CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A5 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A6 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A2 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A6 = CLBLM_L_X8Y118_SLICE_X11Y118_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B3 = CLBLM_R_X11Y116_SLICE_X15Y116_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B4 = CLBLM_L_X12Y119_SLICE_X17Y119_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B5 = CLBLL_L_X4Y120_SLICE_X5Y120_DQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C1 = CLBLM_L_X12Y119_SLICE_X16Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C2 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C3 = CLBLM_L_X10Y120_SLICE_X12Y120_B5Q;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C5 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B5 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D1 = CLBLL_L_X4Y120_SLICE_X5Y120_DQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D2 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D6 = CLBLM_L_X12Y119_SLICE_X17Y119_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D4 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A1 = CLBLM_R_X11Y117_SLICE_X14Y117_DQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A2 = CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A3 = CLBLL_L_X4Y120_SLICE_X5Y120_DQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B1 = CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B3 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_DQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B5 = CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B6 = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C1 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C3 = CLBLM_R_X11Y119_SLICE_X15Y119_B5Q;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C5 = CLBLM_R_X13Y121_SLICE_X18Y121_DQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C6 = CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D2 = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D4 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D5 = CLBLM_R_X11Y121_SLICE_X14Y121_B5Q;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A1 = CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A2 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C1 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A3 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A4 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A6 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A2 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A3 = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A4 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A5 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B6 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C1 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C2 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C4 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C5 = CLBLM_R_X11Y124_SLICE_X14Y124_C5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B2 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B6 = CLBLL_L_X4Y120_SLICE_X4Y120_A5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A4 = CLBLM_L_X12Y119_SLICE_X17Y119_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D1 = CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D2 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D3 = CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D4 = CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C2 = CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B6 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D2 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A1 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A2 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A3 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A4 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A5 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D1 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D2 = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D3 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B4 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B5 = CLBLM_L_X10Y126_SLICE_X12Y126_CO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D4 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D5 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B2 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C4 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A2 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A4 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B2 = CLBLL_L_X4Y120_SLICE_X4Y120_A5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A6 = CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A2 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A3 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B1 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B4 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B5 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C1 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C6 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C1 = CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C2 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C4 = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C5 = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C6 = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D6 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D1 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D3 = CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D1 = CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D2 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D3 = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D4 = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D5 = CLBLL_L_X4Y119_SLICE_X5Y119_DQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D6 = CLBLM_R_X11Y120_SLICE_X15Y120_B5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A2 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A3 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A4 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A5 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B2 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B3 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B4 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B5 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A3 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A5 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A6 = CLBLM_R_X11Y121_SLICE_X15Y121_CQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D1 = CLBLM_R_X11Y124_SLICE_X14Y124_C5Q;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B2 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D2 = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B3 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B4 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B5 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D3 = CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D4 = CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C3 = CLBLM_L_X12Y123_SLICE_X16Y123_DQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C4 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D5 = CLBLM_L_X10Y127_SLICE_X12Y127_DQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A1 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A2 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A3 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D6 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A4 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_A5Q;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D4 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B2 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A3 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A4 = CLBLM_L_X12Y119_SLICE_X16Y119_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A5 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C3 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B5 = CLBLM_R_X11Y120_SLICE_X14Y120_CO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B6 = CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C1 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C3 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C4 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D3 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D2 = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D3 = CLBLM_R_X11Y120_SLICE_X14Y120_DQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D4 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C5 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A1 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_A5Q;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A2 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A3 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A5 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A4 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A3 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B2 = CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B3 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B5 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B1 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B2 = CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C1 = CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C3 = CLBLM_L_X10Y123_SLICE_X12Y123_C5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C6 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A5 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C1 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C3 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A6 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D1 = CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D2 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D3 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D6 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B4 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B6 = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D1 = CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D2 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D3 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D4 = CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A2 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A3 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A1 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D2 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D4 = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B4 = CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B5 = CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B6 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D5 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C1 = CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C3 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C4 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C5 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A2 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A4 = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_AX = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D1 = CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D2 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D3 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C4 = CLBLM_L_X8Y117_SLICE_X10Y117_A5Q;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C5 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C2 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C1 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C2 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C3 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C4 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C6 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D1 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D2 = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D3 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D4 = CLBLL_L_X4Y125_SLICE_X4Y125_AO5;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D5 = CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D2 = CLBLM_L_X8Y116_SLICE_X11Y116_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D3 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D4 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D6 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A2 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A3 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A1 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A2 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A3 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A5 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A6 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B2 = CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B4 = CLBLM_L_X12Y121_SLICE_X16Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B6 = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C2 = CLBLM_R_X11Y121_SLICE_X15Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C3 = CLBLM_R_X11Y122_SLICE_X15Y122_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B2 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C5 = CLBLM_R_X11Y116_SLICE_X15Y116_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D3 = CLBLM_R_X11Y121_SLICE_X15Y121_DQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D4 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B5 = CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D5 = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B6 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A1 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A3 = CLBLM_R_X13Y121_SLICE_X18Y121_DQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A4 = CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B1 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B2 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B5 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C1 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C2 = CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C3 = CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C4 = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C5 = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C2 = CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C6 = CLBLM_L_X10Y121_SLICE_X13Y121_BO5;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C3 = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C4 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D3 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D5 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D6 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A2 = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A4 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A5 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A6 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A1 = CLBLM_R_X11Y124_SLICE_X14Y124_C5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A2 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A4 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A5 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C6 = CLBLM_L_X8Y118_SLICE_X11Y118_CQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D1 = CLBLL_L_X4Y120_SLICE_X5Y120_DQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D2 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B4 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B6 = CLBLM_L_X10Y128_SLICE_X12Y128_AO5;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D3 = CLBLM_L_X10Y118_SLICE_X12Y118_DQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B1 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B3 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B6 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B1 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B2 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D1 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D2 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D3 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D4 = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D5 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D6 = CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A3 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A4 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A5 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B2 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C2 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B3 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B5 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C1 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C2 = CLBLM_R_X11Y122_SLICE_X15Y122_CQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C4 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C3 = CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C5 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C6 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C5 = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C6 = CLBLM_L_X8Y115_SLICE_X11Y115_DQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D1 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D2 = CLBLM_R_X11Y122_SLICE_X15Y122_CQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D3 = CLBLM_R_X11Y122_SLICE_X15Y122_DQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D4 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D5 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A1 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A3 = CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A4 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X25Y143_SLICE_X37Y143_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_AX = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B3 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B4 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A6 = CLBLM_R_X13Y120_SLICE_X19Y120_BO5;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C2 = CLBLM_L_X10Y123_SLICE_X12Y123_DQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C5 = CLBLM_R_X11Y122_SLICE_X14Y122_BO5;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C6 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D1 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D1 = CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D3 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D4 = CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_B5Q;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D3 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D4 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B4 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B5 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C1 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C2 = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C3 = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C4 = CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A5 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C5 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B1 = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B2 = CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C6 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B3 = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B5 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B6 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C3 = CLBLL_L_X4Y120_SLICE_X4Y120_CQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A1 = CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A5 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D1 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D2 = CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B4 = CLBLM_L_X8Y126_SLICE_X11Y126_A5Q;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B6 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C1 = CLBLM_L_X8Y118_SLICE_X11Y118_CQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C2 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C4 = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C6 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D2 = CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D3 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A3 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C1 = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C2 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C3 = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C4 = CLBLM_R_X25Y143_SLICE_X36Y143_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C5 = CLBLM_R_X7Y125_SLICE_X9Y125_DQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C6 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B2 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B5 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C1 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D1 = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D2 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D3 = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D5 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D6 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C4 = CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D1 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D4 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D5 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D6 = CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A2 = CLBLM_R_X11Y122_SLICE_X15Y122_DQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A3 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A4 = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A5 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B2 = CLBLM_L_X12Y122_SLICE_X16Y122_CQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B5 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B6 = CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C2 = CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C4 = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C6 = CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D1 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D5 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D6 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A1 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A2 = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A3 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A4 = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A5 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A6 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B1 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B4 = CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B5 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B6 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C2 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C3 = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C4 = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C6 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D2 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A2 = CLBLM_R_X7Y118_SLICE_X9Y118_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D3 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D4 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D6 = CLBLM_L_X10Y123_SLICE_X12Y123_DQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A5 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A6 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C1 = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B5 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A4 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B4 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C1 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C2 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C4 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C6 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A1 = CLBLM_L_X8Y124_SLICE_X10Y124_A5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D1 = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D2 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D3 = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D4 = CLBLL_L_X4Y127_SLICE_X5Y127_CO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D5 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D6 = CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A6 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A3 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B3 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B6 = CLBLM_R_X11Y124_SLICE_X14Y124_DQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B1 = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B5 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C1 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C2 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C4 = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C6 = CLBLM_L_X8Y122_SLICE_X10Y122_D5Q;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C6 = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D1 = CLBLM_L_X8Y123_SLICE_X11Y123_DQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A1 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A2 = CLBLL_L_X4Y127_SLICE_X5Y127_CO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A3 = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A5 = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A6 = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D2 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A3 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A5 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A6 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B2 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B5 = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C1 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C2 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C3 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D2 = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D3 = CLBLM_L_X10Y119_SLICE_X12Y119_B5Q;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_AX = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B1 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B3 = CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B4 = CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C4 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D1 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D3 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A4 = CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A6 = CLBLM_L_X8Y126_SLICE_X10Y126_A5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B3 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B5 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C2 = CLBLM_R_X11Y124_SLICE_X15Y124_A5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C5 = CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C6 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_L_X12Y117_SLICE_X16Y117_DQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D1 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D2 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D3 = CLBLM_L_X12Y121_SLICE_X16Y121_A5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D4 = CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A1 = CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A2 = CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A3 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A5 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A6 = CLBLM_R_X5Y122_SLICE_X6Y122_A5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B1 = CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B3 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B4 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B5 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B6 = CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D2 = CLBLM_L_X12Y122_SLICE_X16Y122_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A5 = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C2 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C3 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C4 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D5 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D2 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D3 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D4 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A1 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A4 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A5 = CLBLM_L_X8Y123_SLICE_X11Y123_DQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B1 = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B2 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B5 = CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C1 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C2 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C4 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C6 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A1 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A3 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A5 = CLBLL_L_X4Y117_SLICE_X4Y117_C5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A6 = CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D3 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D1 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D2 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A1 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C5 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B2 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B4 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D5 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C1 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C2 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C3 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D1 = CLBLM_L_X8Y121_SLICE_X10Y121_CO5;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D3 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D4 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D5 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D6 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A1 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A2 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A3 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A5 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A6 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B1 = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B2 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B4 = CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B6 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C2 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C3 = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D1 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D3 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D4 = CLBLM_R_X11Y126_SLICE_X15Y126_BO5;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A1 = CLBLM_R_X11Y117_SLICE_X14Y117_DQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A2 = CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A3 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A4 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A5 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B1 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B2 = CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B3 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B4 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B5 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C1 = CLBLM_R_X11Y124_SLICE_X14Y124_C5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C3 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C4 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D1 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D2 = CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D3 = CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D4 = CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D5 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y118_SLICE_X3Y118_A5Q;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B1 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B2 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A3 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A5 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A6 = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B2 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B3 = CLBLM_R_X11Y121_SLICE_X15Y121_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B4 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B5 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C1 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C2 = CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C3 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D2 = CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D5 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C4 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A2 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A3 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A6 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C5 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C6 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B1 = CLBLL_L_X4Y120_SLICE_X5Y120_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B2 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B3 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B4 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C2 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C5 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D3 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A1 = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A2 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A3 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A5 = CLBLM_R_X11Y121_SLICE_X15Y121_DQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A6 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A6 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B1 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B2 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B3 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B4 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B5 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A1 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A2 = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A3 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C1 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C2 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B1 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B2 = CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B5 = CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C2 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D4 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A1 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B5 = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A2 = CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A4 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D1 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D2 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D3 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D4 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D5 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_AX = CLBLM_L_X8Y126_SLICE_X10Y126_A5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B1 = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B2 = CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A1 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A4 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C1 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C2 = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C3 = CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B1 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B4 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B5 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C2 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C3 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C4 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C5 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D2 = CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D3 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D4 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C5 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_SR = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D3 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D5 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D6 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D5 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D4 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D5 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A1 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A6 = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B1 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B2 = CLBLM_L_X8Y123_SLICE_X11Y123_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B4 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B6 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C1 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C2 = CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C3 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C4 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D3 = CLBLM_L_X8Y123_SLICE_X11Y123_DQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D4 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A2 = CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A2 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A3 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A4 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A5 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A5 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B1 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B2 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B3 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B4 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B5 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C2 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C3 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C4 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C5 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B6 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D2 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D3 = CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D4 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D5 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C4 = CLBLM_L_X10Y127_SLICE_X12Y127_DQ;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C5 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A1 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A2 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C6 = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A3 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A4 = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B1 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B2 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B3 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B4 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B5 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B6 = CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A1 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A2 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A5 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C1 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C2 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B1 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B2 = CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B3 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A1 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B4 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B5 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C1 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C6 = CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C3 = CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C5 = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C6 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D4 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A1 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A3 = CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A4 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D2 = CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D3 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A2 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D4 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D6 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A6 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B1 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B3 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A1 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A3 = CLBLM_R_X7Y122_SLICE_X8Y122_B5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A4 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C2 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C3 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B1 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A3 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B5 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D1 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C3 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C4 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C5 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D2 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D3 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D4 = CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D6 = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D1 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D5 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A5 = CLBLM_R_X5Y118_SLICE_X7Y118_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D1 = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C4 = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C5 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A3 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A4 = CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A5 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A6 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D3 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B2 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B5 = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B6 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C3 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C5 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C6 = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D4 = CLBLL_L_X4Y120_SLICE_X4Y120_A5Q;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D4 = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D2 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D3 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D4 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D5 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D5 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D6 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A1 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A2 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A3 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A5 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A6 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_AX = CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B1 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B2 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B3 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B5 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C3 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C4 = CLBLM_L_X10Y119_SLICE_X12Y119_B5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C5 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D6 = CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D3 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D4 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D6 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A5 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B5 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A4 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A5 = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C2 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B2 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B5 = CLBLM_L_X8Y118_SLICE_X11Y118_DO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B6 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D2 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C1 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C2 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C4 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C5 = CLBLM_L_X8Y116_SLICE_X11Y116_CQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C6 = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D2 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D3 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D6 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_AX = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B4 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A1 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A2 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A3 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A4 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A2 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A3 = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B2 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B3 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A4 = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B6 = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A5 = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C3 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A6 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C4 = CLBLL_L_X4Y119_SLICE_X5Y119_CQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D6 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D1 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D2 = CLBLM_R_X7Y118_SLICE_X9Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D3 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D6 = CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B6 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A2 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B2 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A1 = CLBLM_L_X8Y125_SLICE_X11Y125_BO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A3 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A5 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_AX = CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C3 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B2 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B3 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B4 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B5 = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C1 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A2 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A4 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C2 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C4 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A4 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A5 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A6 = CLBLM_R_X7Y125_SLICE_X9Y125_DQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A2 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B2 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B3 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B5 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C1 = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C2 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C3 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C4 = CLBLM_L_X8Y126_SLICE_X11Y126_BO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C5 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D1 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D2 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D4 = CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A3 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D6 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B3 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B5 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C6 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_AX = CLBLM_R_X11Y124_SLICE_X14Y124_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A2 = CLBLM_L_X12Y119_SLICE_X17Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A3 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A4 = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A5 = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_AX = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B4 = CLBLL_L_X4Y120_SLICE_X4Y120_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B5 = CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B6 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_BX = CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C1 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B3 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C2 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C3 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C6 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D1 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D2 = CLBLM_L_X8Y117_SLICE_X10Y117_A5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D4 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D5 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D6 = CLBLL_L_X4Y120_SLICE_X4Y120_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A2 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A5 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B1 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B4 = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B6 = CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C2 = CLBLM_R_X7Y119_SLICE_X9Y119_A5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C3 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C4 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D1 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D2 = CLBLL_L_X4Y119_SLICE_X5Y119_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D3 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D6 = CLBLM_R_X5Y118_SLICE_X7Y118_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D1 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A4 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A5 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D6 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B1 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B2 = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B3 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B4 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B5 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A1 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A4 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A3 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A2 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A4 = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A5 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_AX = CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B2 = CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B3 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B4 = CLBLL_L_X4Y121_SLICE_X5Y121_DQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C1 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C2 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C3 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C4 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C5 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C6 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D1 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D2 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D3 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D6 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X13Y118_SLICE_X19Y118_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A1 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A2 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A3 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A6 = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C2 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B2 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B6 = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C5 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C1 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C2 = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C3 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5 = CLBLL_L_X4Y121_SLICE_X5Y121_DQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C6 = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D2 = CLBLM_L_X8Y126_SLICE_X10Y126_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D4 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D6 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A1 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A2 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A3 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A4 = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A6 = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B1 = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B2 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B4 = CLBLM_L_X8Y125_SLICE_X11Y125_C5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B5 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B6 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C3 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C4 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D2 = CLBLM_R_X5Y124_SLICE_X7Y124_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D3 = CLBLM_L_X8Y125_SLICE_X11Y125_C5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D4 = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5 = CLBLM_L_X8Y122_SLICE_X10Y122_D5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D6 = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A2 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A4 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A5 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A6 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C4 = CLBLM_R_X5Y124_SLICE_X7Y124_A5Q;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C5 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C6 = CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A2 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A4 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A5 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A6 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B2 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B3 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B4 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B5 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B6 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C1 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C2 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C3 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C4 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D1 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D2 = 1'b1;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D1 = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D2 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D3 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D4 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D4 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D5 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A5 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_C5Q;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = CLBLM_R_X7Y118_SLICE_X9Y118_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B4 = CLBLM_L_X8Y126_SLICE_X11Y126_BO5;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B5 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B6 = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C4 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C5 = CLBLM_R_X11Y124_SLICE_X14Y124_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C6 = CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D5 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A1 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A2 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A4 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A5 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B2 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B4 = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B5 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B6 = CLBLM_L_X8Y128_SLICE_X11Y128_AO5;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C1 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C2 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C4 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C5 = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C6 = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D1 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D6 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A2 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A3 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A4 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A6 = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B2 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B3 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B4 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B6 = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C6 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B5 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B3 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C4 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C3 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A1 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A2 = CLBLM_L_X12Y121_SLICE_X16Y121_A5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A3 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A4 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A5 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B2 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B4 = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B5 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C2 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C3 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C4 = CLBLM_L_X8Y122_SLICE_X10Y122_D5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C5 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C5 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D1 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D2 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D3 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D4 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D5 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A1 = CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A6 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B1 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B4 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B5 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C1 = CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C2 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C4 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C5 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D1 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D2 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D3 = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D4 = CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D5 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D6 = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C3 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_L_X12Y117_SLICE_X16Y117_D5Q;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X25Y143_SLICE_X36Y143_AO5;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X25Y143_SLICE_X36Y143_AO5;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A1 = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A2 = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A3 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A4 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A5 = CLBLM_L_X8Y123_SLICE_X11Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A6 = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B1 = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B2 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B3 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B4 = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B5 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B6 = CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C5 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C6 = CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D1 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D2 = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D3 = CLBLL_L_X4Y125_SLICE_X4Y125_AO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D4 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D6 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A1 = CLBLM_L_X12Y123_SLICE_X16Y123_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A2 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A6 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B1 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B2 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B4 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B6 = 1'b1;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C3 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C4 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C5 = CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B1 = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D2 = CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B2 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D4 = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D5 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D3 = CLBLL_L_X4Y125_SLICE_X4Y125_AO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B3 = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B4 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B5 = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C1 = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C2 = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C3 = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C4 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C5 = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C6 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B2 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B3 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D1 = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D6 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D2 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D3 = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A4 = CLBLM_R_X11Y120_SLICE_X14Y120_DQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D4 = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B4 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D5 = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B2 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D6 = CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B5 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B5 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A1 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A2 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A3 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A4 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A5 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B1 = CLBLM_R_X11Y124_SLICE_X15Y124_C5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B2 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B4 = CLBLM_R_X5Y118_SLICE_X7Y118_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B6 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C1 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C2 = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C4 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C5 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C6 = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D2 = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D3 = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D4 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D5 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D6 = CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A1 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A3 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A4 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A5 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B1 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B2 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B3 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B4 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C3 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C4 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C6 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D2 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D4 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D6 = 1'b1;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_L_X12Y117_SLICE_X16Y117_DQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D2 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D3 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D5 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C4 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C5 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A1 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A2 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A3 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A6 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B1 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B2 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B4 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C1 = CLBLM_L_X8Y125_SLICE_X11Y125_C5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C3 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C6 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C4 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C5 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C6 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D1 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D2 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D5 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A2 = CLBLM_R_X3Y120_SLICE_X3Y120_A5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A3 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A4 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A5 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A6 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B2 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B4 = CLBLM_L_X8Y126_SLICE_X10Y126_A5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B5 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B6 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C2 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C3 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_D5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C5 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C6 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_R_X5Y122_SLICE_X6Y122_B5Q;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D2 = CLBLM_R_X11Y126_SLICE_X15Y126_CO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D5 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D6 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X8Y126_SLICE_X11Y126_A5Q;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C4 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C5 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D5 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C5 = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A1 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A2 = CLBLM_R_X5Y118_SLICE_X7Y118_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A3 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A4 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A6 = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B1 = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B2 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B4 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B6 = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C2 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A1 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A2 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C1 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C2 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C3 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D1 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D2 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D3 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D4 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D5 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D6 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D4 = CLBLM_L_X8Y126_SLICE_X10Y126_A5Q;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A3 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A6 = CLBLM_R_X5Y124_SLICE_X7Y124_A5Q;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A1 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A4 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B5 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A1 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A2 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A4 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A6 = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B2 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B4 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B6 = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A1 = CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A2 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A3 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A4 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A5 = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C1 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C2 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C3 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B1 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B2 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B5 = CLBLM_L_X10Y120_SLICE_X12Y120_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D1 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C1 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C2 = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C3 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C4 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D3 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D4 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A4 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D1 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D3 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D4 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A6 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A2 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A3 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A4 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_AX = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B1 = CLBLM_R_X7Y118_SLICE_X9Y118_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B2 = CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B3 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C2 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C3 = CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D2 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D3 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D4 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D5 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A4 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D3 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D4 = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D5 = CLBLM_L_X12Y125_SLICE_X17Y125_BO5;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X7Y122_SLICE_X8Y122_B5Q;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X7Y121_SLICE_X9Y121_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A1 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A2 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A3 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A4 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D6 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A6 = CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B1 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B2 = CLBLM_R_X11Y124_SLICE_X14Y124_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B3 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B4 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B6 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A3 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A4 = CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A5 = CLBLM_L_X12Y118_SLICE_X17Y118_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C3 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B2 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B4 = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B6 = CLBLL_L_X4Y119_SLICE_X5Y119_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C1 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C2 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C4 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B1 = CLBLM_L_X10Y127_SLICE_X12Y127_DQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D2 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D4 = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D6 = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A1 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A2 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A3 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A4 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A5 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B2 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B3 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B5 = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C2 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C5 = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C6 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D2 = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D4 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A1 = CLBLM_R_X13Y118_SLICE_X19Y118_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A4 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B6 = 1'b1;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A4 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B1 = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B2 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B4 = CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B6 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C2 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C3 = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C5 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C6 = CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D1 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D2 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D3 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D4 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D5 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A2 = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A3 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A4 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A6 = CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B1 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B2 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B3 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B4 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B5 = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C3 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C4 = CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D2 = CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D3 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D5 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C4 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C5 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C6 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D6 = CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y118_SLICE_X3Y118_A5Q;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D2 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D3 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A5 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A6 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A2 = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A3 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A6 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C3 = CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B1 = CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B2 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B3 = CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B4 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B6 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C4 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C5 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C1 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C2 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C3 = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C4 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5 = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C6 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D1 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D2 = CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D3 = CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D4 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D6 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B5 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B6 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A2 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A4 = CLBLM_L_X8Y116_SLICE_X11Y116_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B1 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B2 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B6 = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C1 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C2 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C3 = CLBLM_R_X3Y118_SLICE_X3Y118_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D1 = CLBLM_R_X11Y126_SLICE_X15Y126_CO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D2 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D3 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C3 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D2 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D3 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D4 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D5 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D5 = CLBLM_R_X11Y126_SLICE_X15Y126_BO5;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C4 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C5 = CLBLM_L_X12Y123_SLICE_X17Y123_CQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D6 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C6 = CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A5 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A6 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C4 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C6 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B3 = CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B4 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B5 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D2 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C4 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D5 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C5 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C6 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A1 = CLBLM_L_X8Y124_SLICE_X10Y124_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A2 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A3 = CLBLM_R_X5Y122_SLICE_X6Y122_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A4 = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A5 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B1 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B3 = CLBLM_R_X5Y122_SLICE_X6Y122_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B4 = CLBLM_R_X5Y124_SLICE_X7Y124_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B5 = CLBLM_L_X8Y122_SLICE_X10Y122_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B6 = CLBLM_R_X5Y121_SLICE_X7Y121_AO5;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C1 = CLBLM_L_X8Y125_SLICE_X11Y125_C5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C2 = CLBLM_R_X5Y122_SLICE_X6Y122_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C3 = CLBLM_R_X5Y124_SLICE_X7Y124_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C4 = CLBLM_L_X8Y124_SLICE_X10Y124_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C5 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C6 = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D5 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D1 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D3 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D4 = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D5 = CLBLM_L_X8Y122_SLICE_X10Y122_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D6 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A1 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A2 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A3 = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A5 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B2 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B3 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B4 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B5 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C1 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C2 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C3 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C5 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D4 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D6 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_R_X5Y122_SLICE_X6Y122_B5Q;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X13Y118_SLICE_X19Y118_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C5 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A1 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A2 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A3 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A5 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A6 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B1 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B5 = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C1 = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C2 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C3 = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C4 = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C5 = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C6 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D2 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D3 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D4 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D5 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A1 = CLBLM_R_X5Y122_SLICE_X6Y122_B5Q;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A2 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A5 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B3 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B4 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B5 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C2 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C4 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C5 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C6 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D1 = CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D2 = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D3 = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D4 = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D6 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A3 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A5 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A6 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B1 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B2 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B3 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B5 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B6 = CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C2 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C3 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C4 = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D1 = CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D3 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D4 = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D5 = CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D6 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A2 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A6 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B1 = CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B3 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B4 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B6 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C1 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C2 = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C4 = CLBLM_R_X5Y120_SLICE_X6Y120_D5Q;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C5 = CLBLM_R_X25Y143_SLICE_X36Y143_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C6 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D2 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D3 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D4 = CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D5 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D6 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A2 = CLBLM_R_X3Y118_SLICE_X3Y118_A5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A3 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A4 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A6 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B1 = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B2 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B6 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C1 = CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C2 = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C3 = CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C4 = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C5 = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C6 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D1 = CLBLM_L_X10Y124_SLICE_X12Y124_C5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D2 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D4 = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D5 = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D6 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A4 = CLBLM_L_X8Y124_SLICE_X10Y124_A5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A5 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A6 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B1 = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B2 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B4 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B6 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C1 = CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C3 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C4 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C5 = CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C6 = CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D1 = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D2 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D3 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D4 = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D5 = CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D6 = CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B4 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B5 = CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C3 = CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C4 = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C5 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C6 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C2 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D1 = CLBLM_R_X13Y124_SLICE_X19Y124_AO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D2 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D3 = CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C3 = CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D4 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A3 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A5 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B1 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B2 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B3 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B4 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B5 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C3 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C3 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C4 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C6 = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C4 = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C5 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C6 = CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D1 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D3 = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D4 = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D5 = CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D6 = CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B5 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A2 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A4 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A5 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B1 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B2 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B3 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B5 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C1 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_D5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D1 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D2 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D3 = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D4 = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D5 = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D6 = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D3 = CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C2 = CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C3 = CLBLM_R_X13Y125_SLICE_X19Y125_BO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C4 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D5 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C5 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D6 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D5 = CLBLM_R_X13Y126_SLICE_X18Y126_BO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B4 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B5 = CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B6 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C4 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D3 = CLBLM_L_X8Y123_SLICE_X11Y123_DQ;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D6 = CLBLM_L_X10Y123_SLICE_X13Y123_C5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B1 = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B2 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B4 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B5 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B6 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C1 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C2 = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C4 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D1 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D2 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D6 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D5 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A2 = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A3 = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A4 = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A5 = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A6 = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A3 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B2 = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B3 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B4 = CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B5 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B6 = CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C1 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C2 = CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C3 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C4 = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C5 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C6 = CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D2 = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D3 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D4 = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D6 = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B2 = CLBLM_L_X10Y121_SLICE_X13Y121_BO5;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B3 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B4 = CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X25Y143_SLICE_X36Y143_AO5;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X25Y143_SLICE_X36Y143_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A2 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A3 = CLBLL_L_X4Y117_SLICE_X4Y117_C5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A4 = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A6 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B2 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B3 = CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B4 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B5 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A1 = CLBLM_R_X5Y129_SLICE_X6Y129_BO5;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A2 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A4 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B5 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D1 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D2 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D3 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D6 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_AX = CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A1 = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A4 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A5 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_AX = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B1 = CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B4 = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C1 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C3 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D1 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D3 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D4 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D5 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D6 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C6 = 1'b1;
endmodule
