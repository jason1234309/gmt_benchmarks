module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD
  );
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_DO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_DO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AMUX;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BMUX;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_DO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_DO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AMUX;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BMUX;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CMUX;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_AO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_AO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_BO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_BO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_DO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_DO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AMUX;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CMUX;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BMUX;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AMUX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CMUX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d14ff3cdd44ffcc)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_CO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLL_L_X2Y111_SLICE_X1Y111_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fa0a05f5f00ff5f)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_DO6),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3713ff77ff3fffff)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb37fdb77b3ff937f)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb37fb3ffdb3f937f)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a59595999555555)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa33ff33ff)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_DLUT (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbbababafbfbfbba)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_CLUT (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I3(CLBLL_L_X2Y111_SLICE_X0Y111_AO6),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7110fff71000f771)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_DO6),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa55aa563c69c39)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.I3(CLBLL_L_X2Y111_SLICE_X0Y111_AO6),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb4444bbbb4444bb)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_DLUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.I1(CLBLL_L_X2Y112_SLICE_X0Y112_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf0f0b00ffbf0f0b)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_CLUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.I1(CLBLL_L_X2Y112_SLICE_X0Y112_CO6),
.I2(CLBLL_L_X2Y111_SLICE_X0Y111_BO6),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h99cc399c6633c663)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_BO6),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_CO6),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00003f170000ff77)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50f7f7ff75f7ffff)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h20a0b3ff0020a0b3)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.I4(CLBLL_L_X2Y113_SLICE_X0Y113_DO6),
.I5(CLBLL_L_X2Y113_SLICE_X0Y113_BO6),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdbb4af0024b45000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f0ff03c33cc3c)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y113_SLICE_X1Y113_BO6),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CO6),
.I3(CLBLL_L_X2Y113_SLICE_X0Y113_BO6),
.I4(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdb2f4fffcbbf0fff)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b2fbfff3bbfffff)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8727d7d75f5f5f5f)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7888877787777888)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_DO6),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96f05af0a50f96f0)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h043bc4c477884488)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccdfdfa0a05f5f)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X2Y122_SLICE_X0Y122_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(1'b1),
.I4(CLBLL_L_X2Y121_SLICE_X0Y121_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999555500ffffff)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_ALUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_DO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heebbeebb8e2b8822)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_DLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_CO6),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.I4(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.I5(CLBLL_L_X2Y122_SLICE_X0Y122_BO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff153fd5ff40c0)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33c9ff0fcc3600f0)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_CO6),
.I3(CLBLL_L_X2Y122_SLICE_X0Y122_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777788778877)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h020ace460c0c0000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3fcc00cc00)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_ALUT (
.I0(1'b1),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3173717775f7f5ff)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c96963c3c)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3a569f069a53cf0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff66aa9955)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he74d88229a30aa00)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hba4dddff20ffffff)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h317571f573f777ff)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000fff99339933)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0701ff337f1fffff)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd57f2a80b91346ec)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c936c935555ffff)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h137fffff013755ff)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb37f4c80cb0734f8)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a50f0fcc333333)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h03bb2bbb2bff3fff)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5aa5596696699)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d0d4ddd4fdfffff)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbd4d2ddd42b2d222)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0055ff0fff0fff)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff66999999)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bff125abbff22aa)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887887787787788)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7888877787777888)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f053f157f3fff7f)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8e8e8eddeeeeee)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ca0935f935f6ca0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff870fe1c3)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4004d00d0d0d0d0d)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c63f50a39c6f50a)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bbb8eeeafff0aaa)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h59669a55a6666555)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0aafafaf)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9699aa556696aaaa)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dddcfffd444fccc)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936ca05f5fa0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.I4(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h505575f770f7ffff)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I4(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300330033003300)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_CO6),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_CO6),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h28be88eebebeeeee)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h665a9655965a9955)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecb38020fefbc832)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996996666996996)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h60f6c0fcf6f6fcfc)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c96c36996c3693c)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_CO6),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_BO6),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_CO6),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f0fff0fff)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbd422dd24db2dd22)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d4f0ddf4dffddff)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he7654dcf189ab230)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbc433bc4708ff708)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cdf4cdf6c936c93)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdf134cff5f5f00)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3a50f963c5af0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96f0c30f3cf096f0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f7f7f7f7707070)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_BO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5555553333ffff)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h65a69a599a5965a6)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dcfddff8e0ceecc)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he619738c2ad5bf40)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff3f3f3f3f)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he8fa8eafa0e80a8e)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AO6),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_AO6),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_DO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_BO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a959595956a6a6a)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc399699969cc3ccc)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dcfd4fcddff44cc)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbfff3f152a3f00)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_DO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_BO6),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_BO6),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_CO6),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff33ff33ff)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(1'b1),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cc396f0f05a5a)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc33cc3c33c6996)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_CLUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I4(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he8fae8e88eaf8e8e)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c33333ababbbbb)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_ALUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_CO6),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ba459a6f10ef30c)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_CO6),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfaa2a0a2a0fbfa)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_CLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_AO6),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_CO6),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaaa55a65959a6)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_AO6),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_CO6),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f0fff0fff)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1050cf5055000000)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1a3033000f300000)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h14333cccaf003c00)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fd51540ffff3fc0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hac9093a06f90a0a0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd42b2bd4bbbb4444)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_BLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0aaaafff)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_ALUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ac0953f953f6ac0)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h077fffff011f3f3f)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8778ff00e11e33cc)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h222a3bff33bfbfff)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_BLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff5aa5f00f)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88c87f7f7f7fffff)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c6c6c6c93939c6c)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fa0a05f5fff005f)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdfff5f134c5f00)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dcfddffd4fc44cc)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999c33396663ccc)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbd422dd24db2dd22)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8c0fce88e0ccf8e)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a9556a9956aa956)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff77777777)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hed848484ededed84)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd72888777788d728)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h695a96a5a5695a96)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f5f5f5f5f)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf5b271b271a050)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_DLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha66a9a5666aa965a)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_CLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c33c69963cc396)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbd7139f5428ec60a)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_ALUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_CO6),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cccccc39633cc)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c963c963c)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_CO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c63f00f39c6ff00)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AO6),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1073f0ff31f7ffff)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AO6),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c963c963c)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dd4cffcd4d4fcfc)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff999f099f099900)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h63c69c399c3963c6)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff0f0fffff)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3699999693ccccc)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_BLUT (
.I0(CLBLM_L_X8Y119_SLICE_X10Y119_DO6),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_DO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff33ff33ff)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cdfdf4cdfdf4c4c)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he619758a4cb3df20)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdd0d0fdf44040f4)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AO6),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_CO6),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2d22db44b4bb4)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_ALUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AO6),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_CO6),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936ca05f5fa0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_CO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffdf5f135f4c00)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a9696a5a569695a)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_BO6),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_BO6),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AO6),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff0fff0fff)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h27080d0822082208)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h270d484872f24848)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cddc3222dddd222)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcc0cf0cfee0ef0e)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_CLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696669999699966)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f0fff0fff)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0033fff0f0f3ff)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f5f5f5f5f)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(1'b1),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h639cc6399c6339c6)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c96c3693cc3c33c)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcd4f371fcc0f330)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3699999693ccccc)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_DLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8b2c030fcf3e8b2)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_CLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h695aa56996a55a96)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_BLUT (
.I0(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.I1(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff88778877)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7df5ffff14503cf0)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a5aa56996)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_CLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999a55596665aaa)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69963cc3c33c6996)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_ALUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h24046aca2eae6060)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hec75e4f59b571bd7)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h32ddcdddcd223222)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fd51540ffff3fc0)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h93ffc9556c0036aa)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_DLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cc396f0f05a5a)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_CLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996669999666996)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_BLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha05fa05fccdfccdf)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1a1a2200301a2200)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f5f7fff051f557f)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_CLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd788287777d78828)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.I2(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hef8a8aefee8888ee)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a56a9a956)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I1(CLBLM_R_X11Y111_SLICE_X14Y111_AO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_CO6),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h595aa6a5a6a5595a)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_BLUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff33ff33ff)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(1'b1),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h669963cc99999ccc)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1120aa2031200a20)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h06663c3cf6560000)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88778877ffff0077)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h956aa956ff000ff0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.I4(CLBLM_R_X11Y113_SLICE_X15Y113_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699966996699966)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_CLUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.I4(CLBLM_R_X11Y113_SLICE_X15Y113_DO6),
.I5(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf2bf2fb0200b02)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_DO6),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f55ff55ff)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f7f770f770f770)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_DO6),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9cc63c966c36cc66)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999c33396663ccc)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_CO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fcfffff060c66cc)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_CO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h71d4f3fcf550fff0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a956a956a)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_BLUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c3c69c396)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc9396c9c69993ccc)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_BO6),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h456500aa00f00000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a55555ff05ff55)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_ALUT (
.I0(CLBLM_L_X12Y113_SLICE_X16Y113_BO6),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a9696a5a569695a)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_CLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_AO6),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.I4(CLBLM_R_X11Y115_SLICE_X14Y115_CO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0655f30066aa6600)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5f5f5f5f)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf4df4fd0400d04)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_AO6),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.I2(CLBLM_R_X11Y112_SLICE_X14Y112_AO6),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_CO6),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f15bf2abf2abf2a)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_BLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h695a96a5a5695a96)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_ALUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_AO6),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_AO6),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h781e87e187e1781e)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_BO5),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_CO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_AO6),
.I4(CLBLM_R_X11Y115_SLICE_X14Y115_CO6),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_AO6),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ddd8eee8eee8eee)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_DO6),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ca0935f935f6ca0)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_R_X11Y115_SLICE_X14Y115_DO6),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_CO6),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a550fff9a550fff)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_DLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966969999696696)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_AO6),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_CO6),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_BO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_BO5),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_BO6),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0fff0fff)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff00ffffff)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h71d4f3fcf550fff0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33ca55a0ff0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4b44bd22d2dd2)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_AO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_AO6),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_BO6),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f33ff33ff)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd555555ddddffff)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(1'b1),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fffafff06660aaa)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69965aa5a55a6996)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_BO6),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_BO6),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_BO6),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_AO6),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb2dd4ddd4d22b222)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c3963c6c6c6c6c6)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_DLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_BO6),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_DO6),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_DO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff8e8e008e00ff8e)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_AO6),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_AO6),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc333c3335fff0555)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he14b69c378d25af0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he88ea00afaafe88e)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_BO6),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ca0935f935f6ca0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bd4d42bd42b2bd4)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_BO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AO6),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f8fffff07087788)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9aa565a559aaa6aa)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_AO6),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f5555ffff)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c33c69963cc396)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_BO6),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_AO6),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h02ce0c000a460c00)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fb15f93a04ea06c)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0f220ff0f2f02)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h45baba45ba4545ba)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I5(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc333333f0f3f3f3)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f605fa0a05f9f60)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_AO6),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f7f7f780f8f8f8)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969966a55a55aa)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h075570aa8f00da00)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff5f5f5f5f)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_DO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_CO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_BO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff0f0fffff)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_AO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_DO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_CO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_BO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_AO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cccccc3966666)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_DLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_AO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_L_X12Y114_SLICE_X16Y114_AO6),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_DO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaeae00ae00ffae)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_CLUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.I1(CLBLM_L_X12Y112_SLICE_X16Y112_AO6),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_BO6),
.I3(CLBLM_L_X12Y112_SLICE_X16Y112_AO5),
.I4(CLBLM_L_X12Y113_SLICE_X16Y113_BO6),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_CO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h406a705a0af0fa00)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_BO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa9a65aa55659a)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_ALUT (
.I0(CLBLM_L_X12Y113_SLICE_X16Y113_BO6),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_BO6),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_AO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.I4(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.I5(CLBLM_L_X12Y112_SLICE_X16Y112_AO5),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_AO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_DO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_CO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_BO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_AO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a6a6f3f959590c0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_DLUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_L_X12Y114_SLICE_X16Y114_BO6),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_BO6),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_DO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1131aa0a20202020)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_CO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d5530302ea6c0c0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_BO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff007788778877)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y114_SLICE_X16Y114_BO6),
.I4(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_AO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_DO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_CO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_BO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_AO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0bbf2fbfafffffff)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_ALUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haac0960c6ac09ac0)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd42bbbbb2bd44444)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_BLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0223aaff3bbfffff)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_ALUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h575f7fff05570f7f)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9aa65a966a56aa66)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9fa0605f5f9fa060)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c6c936c936c93)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333300000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a95956a6a)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h307077f77377f7ff)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h788778878ff88ff8)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff6c936c93)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b8e8e8ebbeeeeee)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc369693c99cc99cc)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f571f5000a8e0a)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff22bbbbbb)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_DO6),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h57157f377717ff3f)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc66c93c66c6c936c)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h37777fff0307777f)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h95ff6a00a90f56f0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a55a5aaa5aaa5aa)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he9c46ec42508a208)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b8ebbeeaf0affaa)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699cc337711ff33)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_BO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000071f371f371f3)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff69c369c3)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd24b5a0ff05ad24b)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.I4(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2abfbf2abf2abf2a)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ac0953f953f6ac0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f5aa5aa55)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020000000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I2(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_BO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7800ff78ff78ff78)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999a55596665aaa)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h99339933f00f0f0f)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa55555555aaaa)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ffd5fd50554054)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_CO6),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_DO6),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80fe00e8e8ff80fe)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.I2(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3333cc96a55a96)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.I4(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9909660609000600)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6606990906000900)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3693c96693c96c3)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff55ff55ff)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f5f0905ffff9955)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h965a69a566aa9955)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dffddff143c44cc)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f0ff096669996)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b020000bf230000)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_DO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bff02bf02bf002b)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_DO6),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877888777788)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h669696990ff0f00f)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_DO6),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h15ff7fff013357ff)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c93936c6c)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4d2781e3c96f05a)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_BLUT (
.I0(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c30f0faa5500ff)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h93c9cc3c6c36cc3c)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fb3ffff13205fa0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_CO6),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ff70770ff777700)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fa0a05f3f3f3f3f)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.I4(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a959595956a6a6a)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f0f0f00ffffff)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h223f2abf3bbf3fff)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_DO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f07f770f770f770)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f77888877)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3300ff77777777)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h445d5fdf4c5fdfff)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff153fbf3f2a00)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_DO6),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h965aaaaaa59655aa)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a5a6aaaa59a556a)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_DO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee8e8e88dd4d4d44)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_DO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff135fdf5f4c00)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_DO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he26a1d957b3f84c0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f55ff55ff)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h87e1ff33781e00cc)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66aa995573bf8c40)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h550a3ca0390a3ca0)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5500fff0f5f0ff)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999666996669996)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_BO6),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8fce8e88ecf8e8e)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777775f5f5f5f)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc03fc03faabfaabf)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_ALUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h16d0561026e0a6e0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55b9ff13aa4600ec)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h070a0500880aaa00)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he41b7d826c935fa0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_DO6),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h002bbbbb2bffffff)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd52aad527f8007f8)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff69c369c3)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbcd6701acc0c00c0)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0e87f1fff3fffff)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fff7fff077f3f7f)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ca0935f935f6ca0)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h07070f0f01010303)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I3(1'b1),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h577f77ff1537173f)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc69c66966c36cc3c)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5577f7ff77ffffff)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h777fffff173777ff)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c6c935fa0a05f)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69999666a5555aaa)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bbb8eeeafff0aaa)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2db4d24bd24b2db4)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fff030f3cf0c30f)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff55ff55ff)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb42dc3f04bd2c3f0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bb2affab2b2fafa)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a96965a5a)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc369a5a5693cf0f0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f0fff0fff)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(1'b1),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a6a6599a65659a)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966996996996696)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdf134cff5f5f00)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h077fffff011f5f5f)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_CLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4c32df04bc3d2f0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a59955965a66aa)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000100000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bd2b42db42d4bd2)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_CO6),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4d22db44b2dd2)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee8e8e88bb2b2b22)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_BO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a9696a5a569695a)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_CO6),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_CO6),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8eddeecf0cffcc)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4b44bd22d2dd2)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BO6),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1051f3f375f7ffff)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_AO6),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c36c9c936)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he7182bd4639caf50)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_AO6),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff5f5f5f5f)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(1'b1),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cdfdfdf80ececec)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_AO6),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h37077f377f077f7f)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_CO6),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_AO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cf0f0c3960ff0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_BO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h57077f077f577f7f)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_CO6),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_CO6),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8778ff00e11e33cc)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_CO6),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd75f28a0b1934e6c)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_BO6),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_CO6),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6996c3366c6cc6c)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_CO6),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f55ff55ff)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hec80fec880ecc8fe)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_AO6),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_BO6),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_AO6),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdfdfdf134c4c4c)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb44bdd222dd2dd22)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_BO6),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_AO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6639c9c399c9c9c)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_BLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_DO6),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h233b2bff23bfafff)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_ALUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc70fffffe18f3fff)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a59955965a66aa)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_BLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0033ff95959595)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_ALUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h02aa23ff3bffbfff)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6399999639ccccc)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dff143cddff44cc)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hac536f906c935fa0)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22aabbff66aa9955)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffffffffff)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h232b3b3f2fafbfff)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb78877b748778848)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8e71718ef50af50a)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h48de88eededeeeee)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a996655aa)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h639c9c63c63939c6)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f2abf2abf)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h175f0517ffff55ff)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd22d4bb4aa55ff00)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc39969cc69993ccc)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c96c36996c3693c)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff5f5f5f5f)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5f5f5f5f)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8ecf0cddeeffcc)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h93cc6cccc9663666)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h37077f377f077f7f)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5c30f965a3cf0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996696996966996)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_DO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb2cf4d304dcfb230)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4db2b24db24d4db2)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_DO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bffbbff125a22aa)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(CLBLM_R_X11Y114_SLICE_X15Y114_CO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff55ff55ff)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f60c03f3fc09f60)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_DO6),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc369a5a5693cf0f0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h03af2baf2bff3fff)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_DO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a6a6599a65659a)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff77777777)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb478d21e3cf0965a)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696969999696966)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I2(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc69963cc39999ccc)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f3f3f3f3f)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96996696cc33cccc)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_CO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf999fff990009990)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_CO6),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_CO6),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c6c6399c63639c)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_CO6),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_CO6),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.I5(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff0fff0fff)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dddd444cffffccc)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h10f531f573fff7ff)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_CLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_BLUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5965a965a965a)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ff70770f7f77070)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_DO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_BO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbfff3f152a3f00)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hec80b320fec8fb32)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_DLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_AO5),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_BO6),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c36c9c936)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_CLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_AO5),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_BO6),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h965aaaaaa59655aa)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0fff0fff)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9999000fff99990)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_DLUT (
.I0(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_AO6),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966666699996)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_CLUT (
.I0(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_AO6),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_DO6),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff0f0fffff)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(1'b1),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4d22db44b2dd2)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_AO6),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_DO6),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_BO6),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c96c36996c3693c)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_BLUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_CO6),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_DO6),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_DO6),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0fff0fff)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5070757777f7f7ff)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_DO6),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc96c399c693c99cc)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_BLUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc96c693c399c99cc)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_DO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f07f770ff777700)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877888777788)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996996696966666)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h659a9a65a65959a6)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_BO6),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AO6),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_CO6),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hef8aae08df455d04)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_BO6),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h659aa6599a6559a6)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_BO6),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h95ff6a00a93356cc)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_BO6),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777773f3f3f3f)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a956a957b843fc0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee8888eefec8c8fe)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha66599aa599a99aa)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_AO5),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_AO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0df2f20df20d0df2)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ff70770f7f77070)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_CO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969699666666)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_CO6),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f5555ffff)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h93c9cc666c36cc66)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_DLUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_AO6),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0320f02023205020)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h345834a84458b4a8)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88778877ffff0077)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff5f5f5f5f)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf11101c10505ffff)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c9ca0606c6ca0a0)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a4bbbbba5b44444)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_BLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0baaffafbfffff)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_ALUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fffffffff)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha66a66aa9955a66a)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_DLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaafb22bb22ba00a)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_CLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I4(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c3c69c396)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_BLUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff5f5f5f5f)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff55ff55ff)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_DO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_CO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_BO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h695a96a5a5695a96)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_CO6),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_AO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_BO6),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_CO6),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_AO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_CO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_BO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_AO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999999659aaaaa)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_BO6),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcc0f330fec8fb32)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_AO5),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_BO6),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h693c696996c39696)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_BO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_AO5),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff3f3f3f3f)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bf3ffff12305af0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_CO6),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33ca55a0ff0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h48dedede88eeeeee)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_BLUT (
.I0(CLBLM_L_X12Y113_SLICE_X16Y113_DO6),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c996633cc)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c3f05a3c96f05a)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_R_X11Y112_SLICE_X14Y112_AO6),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f5d450f3fffcf0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_DO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_L_X12Y114_SLICE_X16Y114_DO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c3693c993c96c36)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_BLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_DO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_BO6),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_AO6),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_AO6),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_CO6),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777775f5f5f5f)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd25a78f0b4961e3c)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_CO6),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_BO6),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1322b1000022aa00)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777733ff33ff)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha699599965aa9aaa)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_DLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_R_X11Y115_SLICE_X14Y115_BO6),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9909090f9f9f990)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_CLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_AO6),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.I5(CLBLM_R_X11Y115_SLICE_X14Y115_BO6),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a95956a6a)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_BLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_L_X12Y114_SLICE_X16Y114_DO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c3693c993c96c36)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_BO6),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_AO6),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb2cf4dcf4d30b230)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_AO5),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_AO5),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X12Y114_SLICE_X16Y114_DO6),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936ca05f5fa0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h48de88eededeeeee)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_BLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c6c93936c6c9c6c)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_DO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96669996cccc3c3c)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_R_X11Y116_SLICE_X15Y116_CO6),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hecb38020fefbc832)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.I1(CLBLM_R_X11Y116_SLICE_X15Y116_CO6),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AO5),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_BO6),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a9696a5a569695a)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AO5),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_BO6),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_CO6),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f33ff33ff)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccff33ce083b02)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_DLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_AO6),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_BO6),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_AO5),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_AO6),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_BO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c3c69c396)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_AO6),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_AO6),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_AO6),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_DO6),
.I5(CLBLM_R_X11Y116_SLICE_X15Y116_BO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696669999699966)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_BLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_AO6),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_BO6),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_BO6),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_AO6),
.I5(CLBLM_R_X11Y116_SLICE_X15Y116_AO5),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff5f5f5f5f)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ff7ff7707707700)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cccccc6963666)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_CLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_BO6),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877888777788)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h036cf060636c5060)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f7f770f770f770)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c3c6cccc6963666)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_CLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_AO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999c33396663ccc)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_CO6),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000fffcccccfff)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(1'b0),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X1Y112_DO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X1Y112_BO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_CO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_AMUX = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_AMUX = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_BMUX = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_CMUX = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_DMUX = CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_AMUX = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_AMUX = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_AMUX = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_BMUX = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_CMUX = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_AMUX = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_AMUX = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_AMUX = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_CMUX = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_AMUX = CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_BMUX = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_CMUX = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_AMUX = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_AMUX = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_AMUX = CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_AMUX = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_BMUX = CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_AMUX = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_AMUX = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_CMUX = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_AMUX = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_BMUX = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_BMUX = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_AMUX = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_AMUX = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_AMUX = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_AMUX = CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_BMUX = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_AMUX = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_BMUX = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_CMUX = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A = CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_AMUX = CLBLL_L_X4Y121_SLICE_X4Y121_AO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A = CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_AMUX = CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A = CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_AMUX = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_CMUX = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_AMUX = CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_CMUX = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_AMUX = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_AMUX = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_DMUX = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_AMUX = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_DMUX = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_AMUX = CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_AMUX = CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A = CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B = CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C = CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A = CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_AMUX = CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C = CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_AMUX = CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A = CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_AMUX = CLBLM_L_X8Y121_SLICE_X11Y121_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_CMUX = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_AMUX = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_AMUX = CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_DMUX = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_AMUX = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_AMUX = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_BMUX = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_CMUX = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_AMUX = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_BMUX = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_AMUX = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_AMUX = CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_AMUX = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B = CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C = CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D = CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_AMUX = CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A = CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B = CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_AMUX = CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_BMUX = CLBLM_L_X10Y116_SLICE_X12Y116_BO5;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A = CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_AMUX = CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A = CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_AMUX = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_CMUX = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_BMUX = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_AMUX = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_AMUX = CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_CMUX = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_AMUX = CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A = CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B = CLBLM_L_X12Y112_SLICE_X16Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C = CLBLM_L_X12Y112_SLICE_X16Y112_CO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D = CLBLM_L_X12Y112_SLICE_X16Y112_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_AMUX = CLBLM_L_X12Y112_SLICE_X16Y112_AO5;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A = CLBLM_L_X12Y112_SLICE_X17Y112_AO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B = CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C = CLBLM_L_X12Y112_SLICE_X17Y112_CO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A = CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C = CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D = CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_AMUX = CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_BMUX = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A = CLBLM_L_X12Y113_SLICE_X17Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B = CLBLM_L_X12Y113_SLICE_X17Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C = CLBLM_L_X12Y113_SLICE_X17Y113_CO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D = CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A = CLBLM_L_X12Y114_SLICE_X16Y114_AO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_AMUX = CLBLM_L_X12Y114_SLICE_X16Y114_AO5;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_BMUX = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_CMUX = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A = CLBLM_L_X12Y114_SLICE_X17Y114_AO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B = CLBLM_L_X12Y114_SLICE_X17Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C = CLBLM_L_X12Y114_SLICE_X17Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D = CLBLM_L_X12Y114_SLICE_X17Y114_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_AMUX = CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_CMUX = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AMUX = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_AMUX = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_AMUX = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_AMUX = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AMUX = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_BMUX = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_AMUX = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_AMUX = CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_AMUX = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_BMUX = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_CMUX = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_AMUX = CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_AMUX = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_CMUX = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_DMUX = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_AMUX = CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_AMUX = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_AMUX = CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_CMUX = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_AMUX = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_AMUX = CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_BMUX = CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_CMUX = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_AMUX = CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_AMUX = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_DMUX = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_AMUX = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_BMUX = CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_AMUX = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_AMUX = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_DMUX = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_AMUX = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_AMUX = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_AMUX = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_CMUX = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_AMUX = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_BMUX = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_BMUX = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_AMUX = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CMUX = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_BMUX = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_AMUX = CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_AMUX = CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_AMUX = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_CMUX = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_AMUX = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_CMUX = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_AMUX = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_BMUX = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_AMUX = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_BMUX = CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_AMUX = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_AMUX = CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_AMUX = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_AMUX = CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_BMUX = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_BMUX = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_CMUX = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B = CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_AMUX = CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_AMUX = CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_DMUX = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_AMUX = CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_BMUX = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_AMUX = CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_DMUX = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_AMUX = CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_AMUX = CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_CMUX = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A = CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_AMUX = CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_AMUX = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_AMUX = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_AMUX = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_AMUX = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C = CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D = CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A = CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_AMUX = CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_DMUX = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B = CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_AMUX = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D = CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_AMUX = CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_DMUX = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A = CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_AMUX = CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_AMUX = CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_CMUX = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_AMUX = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_CMUX = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A = CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_AMUX = CLBLM_R_X11Y117_SLICE_X15Y117_AO5;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A2 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A3 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A4 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B2 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B3 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B4 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C2 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C3 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C4 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D2 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D3 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D4 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A3 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A4 = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A5 = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D5 = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D6 = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A1 = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A4 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C4 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C5 = CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C6 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D1 = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D2 = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D3 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D4 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D5 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D6 = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A3 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A4 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C5 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C6 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D2 = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D6 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B2 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B4 = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B6 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C3 = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D3 = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D4 = CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D4 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A3 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A4 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B1 = CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B2 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B3 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B4 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B5 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B6 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C2 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C1 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C2 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C3 = CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C4 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C5 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C6 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C5 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D1 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D2 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D6 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A1 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A2 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A3 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A4 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A5 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A6 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B1 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B2 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B3 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B4 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B5 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B6 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C1 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C2 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C3 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C4 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C5 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C6 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D2 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D4 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D5 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D6 = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A4 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A5 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B1 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B2 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B6 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A1 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A2 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A3 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A4 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A5 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A6 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B1 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B6 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C1 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C2 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C3 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C4 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C5 = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C6 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D3 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D6 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A2 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A3 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B4 = CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B5 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C1 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C4 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C6 = CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A2 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A4 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A5 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B1 = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B2 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B3 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B4 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B5 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B6 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C1 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C3 = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C5 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D1 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D5 = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D6 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A3 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A4 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A5 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D1 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D2 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D5 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A1 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A3 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B1 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B2 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B3 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B4 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B5 = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B6 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C1 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C2 = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C4 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C5 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C6 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D1 = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D2 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D3 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D4 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D5 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D6 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A2 = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A6 = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B2 = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B6 = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C1 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C4 = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D3 = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D4 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A2 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B1 = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B2 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B3 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B4 = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B5 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B6 = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C1 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C2 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C3 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C4 = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C5 = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C6 = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D3 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D4 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D5 = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A1 = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A4 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C1 = CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C2 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C5 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D4 = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D6 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A1 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A2 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A3 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A4 = CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A5 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A6 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B1 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B4 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C3 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C4 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A1 = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A2 = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A3 = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A4 = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A5 = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A6 = CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B1 = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B4 = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C3 = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C4 = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D1 = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D2 = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D3 = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D4 = CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D5 = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D6 = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C3 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C1 = CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C6 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D6 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A6 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B5 = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B6 = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C1 = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C2 = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D2 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D3 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D4 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B6 = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = 1'b0;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A1 = CLBLM_L_X10Y116_SLICE_X12Y116_BO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A2 = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A3 = CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A4 = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A5 = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A6 = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B2 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B3 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B4 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C2 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C3 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C4 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D2 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D3 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D4 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A1 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A4 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A6 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B1 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B2 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B6 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A5 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A6 = 1'b1;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B1 = CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B2 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B3 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B4 = CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B5 = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B6 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C4 = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D3 = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D4 = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A2 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B2 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C1 = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C2 = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C4 = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_BO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C4 = CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B1 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B2 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B3 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B4 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B5 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B6 = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C1 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C2 = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C4 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C5 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C6 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D1 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D5 = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D6 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A2 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A5 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B2 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B3 = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B4 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B5 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C1 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C2 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C4 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C5 = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C6 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D1 = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D2 = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A2 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A6 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B5 = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B6 = CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B4 = CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C1 = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C6 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C4 = CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C5 = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B4 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A5 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A6 = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C1 = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D6 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A2 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A3 = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A4 = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A6 = CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B5 = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B6 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C2 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C6 = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C4 = CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C5 = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A5 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B1 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B2 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B5 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C2 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D4 = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D5 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C6 = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B3 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B5 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C3 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C5 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D3 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D5 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A1 = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A2 = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A3 = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A4 = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A5 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A6 = CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B3 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B5 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C3 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C5 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D3 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D5 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A2 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A3 = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B1 = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B2 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B3 = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B4 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B5 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B6 = CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C4 = CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A4 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C6 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A5 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C1 = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C2 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C3 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B2 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D2 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D4 = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D6 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B5 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B6 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B1 = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B2 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B3 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B5 = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B6 = CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C2 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C3 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A3 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A4 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B5 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B6 = CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C2 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C4 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C6 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D2 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D3 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D6 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A2 = CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B1 = CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B2 = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C3 = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C4 = CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D6 = CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B1 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B2 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B3 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B4 = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B6 = CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C3 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C5 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C6 = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D1 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D2 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D6 = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D4 = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D5 = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D6 = CLBLM_L_X8Y121_SLICE_X11Y121_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C2 = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C3 = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C6 = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B1 = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B3 = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B4 = CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B5 = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B6 = CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C3 = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C5 = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D1 = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D3 = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D4 = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A2 = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A5 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A6 = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B1 = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C4 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C5 = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D2 = CLBLM_R_X11Y117_SLICE_X15Y117_AO5;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D3 = CLBLM_L_X12Y114_SLICE_X16Y114_AO5;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D6 = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A1 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A2 = CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A3 = CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A4 = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A5 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A6 = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B1 = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B5 = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C1 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C2 = CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C3 = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C4 = CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C5 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C6 = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D2 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D6 = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B1 = CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B2 = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B3 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B4 = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B5 = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B6 = CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C1 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C2 = CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C3 = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C4 = CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C5 = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C6 = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D1 = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D2 = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D3 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D4 = CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D5 = CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D6 = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B3 = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B4 = CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B5 = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B6 = CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C1 = CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C2 = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C3 = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C4 = CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C6 = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D2 = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D3 = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D5 = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A2 = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A5 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B6 = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C1 = CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C2 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D3 = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D4 = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B4 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B5 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C1 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C2 = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C6 = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D4 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D6 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A1 = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A3 = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A6 = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B1 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B3 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B4 = CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B5 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B6 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C3 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C5 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C1 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D1 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D2 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D3 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D5 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D6 = CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A1 = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A5 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B1 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B6 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C6 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A1 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A3 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A4 = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B1 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B2 = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B3 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A1 = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A2 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A4 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A2 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A3 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B2 = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B3 = CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B4 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C1 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B5 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B6 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C4 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C2 = CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C6 = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C3 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C5 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B2 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B3 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C2 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D1 = CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D3 = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D5 = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D2 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A3 = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A4 = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A6 = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B4 = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B6 = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A1 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C2 = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C3 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B1 = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B2 = CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B3 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C2 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B5 = CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C5 = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C6 = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C1 = CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D4 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D6 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D2 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D3 = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D4 = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D3 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D4 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A3 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A4 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B1 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B2 = CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B4 = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B6 = CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B3 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C1 = CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C3 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B3 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C5 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C3 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C4 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D4 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D3 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A5 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B1 = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B2 = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A1 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A2 = CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A3 = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A4 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A5 = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A6 = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A4 = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B1 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B4 = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B6 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B5 = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B6 = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C2 = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C4 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C2 = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C4 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C5 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D2 = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D5 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A1 = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A2 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A3 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A6 = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B6 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C5 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D4 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A1 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A1 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A2 = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A3 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A4 = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A5 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B1 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B2 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B3 = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B4 = CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B5 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B6 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B1 = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B2 = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C1 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C2 = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C3 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C4 = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C5 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C6 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B5 = CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B6 = CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C5 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D1 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D5 = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D4 = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D5 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A1 = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A2 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A4 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A5 = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B1 = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B2 = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B3 = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B4 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B5 = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B6 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C1 = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C2 = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C3 = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C5 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C6 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D1 = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D2 = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D4 = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D5 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A3 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A5 = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B2 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B4 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C2 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C4 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D2 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D4 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B1 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B2 = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B4 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B3 = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C1 = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C2 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C3 = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C4 = CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C5 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C6 = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D1 = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D2 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D5 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B1 = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B3 = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B4 = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B5 = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B6 = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C1 = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C2 = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C3 = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C4 = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C5 = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D2 = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D4 = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D5 = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B1 = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B2 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B5 = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C1 = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C2 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C3 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C4 = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C5 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D3 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D5 = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B2 = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B3 = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B2 = CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B3 = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B4 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A2 = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A6 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B4 = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B6 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C5 = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D3 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A1 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A3 = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B1 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B2 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B4 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B6 = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C1 = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C3 = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C6 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D2 = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D5 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A2 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A6 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B2 = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B6 = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A5 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A6 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C1 = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C2 = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C3 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B6 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D1 = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D2 = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C4 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D3 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D4 = CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A2 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D4 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B4 = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A2 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A3 = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A6 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C1 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C2 = CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C3 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B3 = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B4 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B5 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D1 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D2 = CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D3 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C2 = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C6 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D4 = CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D6 = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D2 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D4 = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D5 = CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B1 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A1 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A2 = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A4 = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B1 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B2 = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C3 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B1 = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B2 = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B3 = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B4 = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B5 = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C2 = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B2 = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5 = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B6 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C4 = CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5 = CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C6 = CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C2 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5 = CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D6 = CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D2 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A1 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A2 = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A3 = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A4 = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A6 = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B1 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C4 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C3 = CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A1 = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = CLBLL_L_X4Y121_SLICE_X4Y121_AO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D2 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D3 = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D6 = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B3 = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B4 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C6 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A4 = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A5 = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D1 = CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D2 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D4 = CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A1 = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B2 = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B5 = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D3 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D5 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D6 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A4 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B3 = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B4 = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B6 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C5 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C6 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D1 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D2 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D3 = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D4 = CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D5 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D6 = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C4 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A1 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A2 = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A3 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A4 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A5 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A6 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B1 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B2 = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B3 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B6 = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C2 = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C3 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C4 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C5 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A1 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A6 = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B3 = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B5 = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C1 = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C3 = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C6 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D4 = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D5 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C5 = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D3 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B5 = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B6 = CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C3 = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A1 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A4 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A6 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B1 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B2 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B6 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C5 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A3 = CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A6 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B6 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B4 = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A1 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D2 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D6 = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A2 = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A5 = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A6 = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B2 = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B4 = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B6 = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C4 = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C6 = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B2 = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B4 = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C2 = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D1 = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D2 = CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D6 = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B2 = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B1 = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B4 = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C3 = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C6 = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C4 = CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C5 = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C6 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOB33_X0Y133_IOB_X0Y134_O = 1'b0;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D5 = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D6 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C6 = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B6 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D3 = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D4 = CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C4 = CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5 = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C6 = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B4 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C4 = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C6 = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A4 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A6 = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B3 = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B4 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A3 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A4 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B1 = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B3 = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B4 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C2 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C5 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D2 = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D5 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D6 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A4 = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A5 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B1 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B2 = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C5 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C5 = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C6 = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A1 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A3 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A4 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A5 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B1 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B3 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B4 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B5 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C1 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C3 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C4 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C5 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D1 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D3 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D4 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D5 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A1 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D3 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B1 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B3 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B4 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B5 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C1 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C4 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C5 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D1 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D3 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D4 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D5 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B6 = CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C5 = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C6 = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A1 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A3 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A5 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B1 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B3 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B5 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C1 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C3 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C5 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D1 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D3 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D5 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A1 = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A2 = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A3 = CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A4 = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A5 = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A6 = CLBLM_L_X12Y112_SLICE_X16Y112_AO5;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C1 = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C2 = CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C3 = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C4 = CLBLM_L_X12Y112_SLICE_X16Y112_AO5;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C5 = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C6 = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D1 = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D6 = CLBLM_L_X12Y114_SLICE_X16Y114_AO6;
endmodule
