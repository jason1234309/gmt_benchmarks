module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y119_IOB_X0Y119_IPAD,
  input LIOB33_X0Y119_IOB_X0Y120_IPAD,
  input LIOB33_X0Y121_IOB_X0Y121_IPAD,
  input LIOB33_X0Y121_IOB_X0Y122_IPAD,
  input LIOB33_X0Y123_IOB_X0Y123_IPAD,
  input LIOB33_X0Y123_IOB_X0Y124_IPAD,
  input LIOB33_X0Y125_IOB_X0Y125_IPAD,
  input LIOB33_X0Y125_IOB_X0Y126_IPAD,
  input LIOB33_X0Y127_IOB_X0Y127_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD
  );
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AMUX;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AMUX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AMUX;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_BO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_CO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_DO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_BO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_BO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_CO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_CO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_DO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AMUX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffafffaff)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(1'b1),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(1'b1),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeeffffffff)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(1'b1),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbfbfbfffffffb)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(CLBLL_L_X2Y113_SLICE_X0Y113_DO6),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff3fff2ff)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLL_L_X2Y113_SLICE_X0Y113_CO6),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88008800dd00dd00)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h75307530ffffffff)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f01100000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.I5(CLBLL_L_X2Y113_SLICE_X1Y113_CO6),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f5f3f0f77553300)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffff7fffff)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000400040404000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_BO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5510551055005500)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_DLUT (
.I0(CLBLL_L_X2Y116_SLICE_X0Y116_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0f5f5f57035757)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_CLUT (
.I0(CLBLL_L_X2Y113_SLICE_X0Y113_AO6),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_DO6),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLL_L_X2Y116_SLICE_X0Y116_BO6),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0203030300030303)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33100100af000500)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y127_IOB_X0Y127_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffbf00ffff)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.I3(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff44ff04)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_BO6),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I5(CLBLL_L_X2Y116_SLICE_X1Y116_CO6),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808000000880000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafafa88aaf8fa)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_DLUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(LIOB33_X0Y125_IOB_X0Y125_I),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y123_IOB_X0Y124_I),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffbffffff)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y119_IOB_X0Y120_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000101e8e88080)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(1'b1),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44cc44cceefffafa)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff0055000f0007)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_DLUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I3(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_DO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_CLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_BLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I4(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I5(CLBLL_L_X2Y117_SLICE_X1Y117_CO6),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffefffefffff)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_ALUT (
.I0(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c5c5c5c5c5f5c5f)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_CLUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(1'b1),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y119_IOB_X0Y120_I),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002245cd45cd)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0e0f0f0f)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_DLUT (
.I0(LIOB33_X0Y123_IOB_X0Y124_I),
.I1(LIOB33_X0Y125_IOB_X0Y125_I),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I3(LIOB33_X0Y123_IOB_X0Y123_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(CLBLL_L_X2Y117_SLICE_X0Y117_BO6),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000100010000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_CLUT (
.I0(CLBLL_L_X2Y116_SLICE_X1Y116_AO5),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_BO6),
.I3(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00330033bbffaaaa)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_BLUT (
.I0(CLBLL_L_X2Y116_SLICE_X0Y116_DO6),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(1'b1),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003370730000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(LIOB33_X0Y121_IOB_X0Y121_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h575703035f5f0303)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_CLUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(1'b1),
.I4(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I5(CLBLL_L_X2Y117_SLICE_X0Y117_BO6),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffbfff)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y119_IOB_X0Y120_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeff4ef000ffff)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y127_IOB_X0Y127_I),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777777777777)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a0a0a0a08)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffbbbf)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_BLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05ff05ffcc008000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cfffff55df55df)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.I3(CLBLL_L_X2Y116_SLICE_X1Y116_BO6),
.I4(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00050004000400)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y125_IOB_X0Y125_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(LIOB33_X0Y123_IOB_X0Y124_I),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcfdf0000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I1(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_DO6),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc0ccbbbbbfbb)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y121_IOB_X0Y121_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33133313ffffffff)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001030)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I5(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcaaaaffccaaaa)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I4(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000a80000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.I3(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050ffff505cffff)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I2(CLBLL_L_X2Y116_SLICE_X0Y116_DO6),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h03ff030300a80000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_ALUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff30303030)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0e0e0e0e0e0f0f)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_CLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I3(1'b1),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5c0d5f0f0c0c0)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_BLUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I1(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h337f337fa0a0a0a0)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha00a820a0a0a0a0a)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_DLUT (
.I0(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffee0000afae)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_CLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f1fff0f0ffff)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I4(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cc00ff03ff03)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaafaaafafafae)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_DLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I3(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdffffffff)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_CLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_DO6),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_CO6),
.I3(CLBLL_L_X2Y122_SLICE_X0Y122_DO6),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_DO6),
.I5(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f1f500000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_BLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff55550010)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_ALUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffca880008000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_ALUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaabaaaa)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_CLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.I1(CLBLL_L_X2Y122_SLICE_X0Y122_CO6),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I3(CLBLL_L_X2Y122_SLICE_X0Y122_DO6),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_CO6),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefffff)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I1(CLBLL_L_X2Y122_SLICE_X0Y122_CO6),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_CO6),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.I5(CLBLL_L_X2Y122_SLICE_X0Y122_DO6),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000ff00ff)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I1(CLBLL_L_X2Y122_SLICE_X0Y122_CO6),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_CO6),
.I4(CLBLL_L_X2Y122_SLICE_X0Y122_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_DO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_CO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_BO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_DO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_CO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_BO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffffffefefefef)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfffffffeff)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(LIOB33_X0Y123_IOB_X0Y124_I),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff55555554)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(LIOB33_X0Y123_IOB_X0Y124_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3fffffaa2aaaaa)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(LIOB33_X0Y123_IOB_X0Y123_I),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000011f0f0f0e0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccfcffff)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y123_IOB_X0Y123_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8fafafafafafafa)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffe8aaaaaaa)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(LIOB33_X0Y123_IOB_X0Y123_I),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0faaaaffffffff)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(1'b1),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f333f332f222f22)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I3(LIOB33_X0Y123_IOB_X0Y123_I),
.I4(1'b1),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4400000005050505)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I1(LIOB33_X0Y123_IOB_X0Y124_I),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbfbfbfae)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_CO6),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8808aa0acc0cff0f)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff00fffffe30)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0c080f0f0c0c0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(CLBLL_L_X4Y116_SLICE_X5Y116_BO6),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_CO6),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0444000000000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b8fffff8b888b88)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y123_IOB_X0Y123_I),
.I5(LIOB33_X0Y123_IOB_X0Y124_I),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a0030002a002a2a)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30300000ff45ff55)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003300330033)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h003700ffc8c80000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222220000aa0088)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y119_IOB_X0Y120_I),
.I2(1'b1),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y121_IOB_X0Y121_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h23220002a0aa000a)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff22ff2022222020)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y121_IOB_X0Y121_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h005000500000cecc)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(LIOB33_X0Y123_IOB_X0Y124_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h550055005500ffff)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y119_IOB_X1Y120_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaabaabaaabbaa)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(RIOB33_X105Y119_IOB_X1Y120_I),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7020002070770000)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(LIOB33_X0Y123_IOB_X0Y123_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafca0fcaa00a000)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y121_IOB_X0Y121_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0fff0f3f0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_DO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aff0ace0fff0fcf)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33f300000f0f)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffeeffefefeeee)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3b3bfbfb)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(1'b1),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3bffff3f3b3f3b)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff7fff75)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(LIOB33_X0Y127_IOB_X0Y127_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3fff2fffffffe)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0300000a02)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.I5(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecccecccccccecc)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.I1(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30000000a0a0a2a0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffce33333131)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_X0Y127_IOB_X0Y127_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0b00000b0b000bb)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I1(LIOB33_X0Y123_IOB_X0Y124_I),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hceffffffceffceff)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3303bbab)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_DO6),
.I1(CLBLL_L_X2Y113_SLICE_X0Y113_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0d0d0dd00000000)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0700000f0200000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaaaaab)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe8ff8000000000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c5c5f5f00000202)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(1'b1),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000000000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_DLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3322322222222222)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbbaabfaf)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.I2(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.I3(CLBLL_L_X2Y118_SLICE_X1Y118_AO6),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000f30000000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050f0f0f0f0f0f0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd55ffffd050f0f0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f111111ff111111)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_BLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333303030303030)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee88ee8888008800)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a0a0a000aaa0aa)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(1'b1),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y121_IOB_X0Y121_I),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000055fd)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_BLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.I5(CLBLL_L_X2Y117_SLICE_X1Y117_DO6),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444545444ff54ff)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(LIOB33_X0Y123_IOB_X0Y123_I),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffddffcc0f0c)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.I1(CLBLL_L_X2Y116_SLICE_X0Y116_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_CO6),
.I4(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11111111ffff1f11)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0eacfefc0eaeaea)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y127_IOB_X0Y127_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h300000000fffffff)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7070000070705050)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(1'b1),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(LIOB33_X0Y121_IOB_X0Y121_I),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000000)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y119_IOB_X0Y120_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000504)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0000000eaaaaaaa)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I1(RIOB33_X105Y119_IOB_X1Y120_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444044ccccc0cc)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_DO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7530303030303030)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I1(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004aaae0044aaee)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(CLBLL_L_X2Y116_SLICE_X0Y116_DO6),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fe0000000101)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd0000dd000000)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I2(1'b1),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_DO6),
.I5(RIOB33_X105Y119_IOB_X1Y120_I),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdc0050505000)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.I4(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ccc0fff08880aaa)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00a000880080)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I1(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.I2(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc00000008)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff30ff31ffffffff)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303030303031)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff85ff80)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000feeef000f)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(LIOB33_X0Y119_IOB_X0Y120_I),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303030003030301)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(RIOB33_X105Y119_IOB_X1Y119_I),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_DO6),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_DO6),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeae0000aeff0000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf8fffaf0f0f0f0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.I4(RIOB33_X105Y119_IOB_X1Y120_I),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020002000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_DLUT (
.I0(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888d8d8d8c)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_CLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333337f7f7f)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc80cccc8080)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fc00fc00a800a8)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.I2(LIOB33_X0Y127_IOB_X0Y127_I),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.I4(1'b1),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffcc0000f0c0)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c840000000cc)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_BLUT (
.I0(CLBLL_L_X2Y116_SLICE_X0Y116_DO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaab00000003)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_ALUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fe54fe54)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_DLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I3(CLBLM_R_X3Y123_SLICE_X2Y123_AO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0000000f00010)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_CLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_DO6),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff55555554)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_BLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_DO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfe00000000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000888a)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_CLUT (
.I0(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333200000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5455445550550055)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_ALUT (
.I0(CLBLL_L_X2Y116_SLICE_X0Y116_DO6),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddddddffddff)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I2(1'b1),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(1'b1),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y119_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y119_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y120_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y120_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y121_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y121_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y122_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y124_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y125_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y126_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y127_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X2Y123_SLICE_X0Y123_AO5),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X0Y118_CO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLL_L_X2Y123_SLICE_X0Y123_AO6),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_CO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_BO6),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_DO6),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X0Y122_BO6),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLL_L_X2Y125_SLICE_X0Y125_BO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X2Y125_SLICE_X0Y125_AO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLL_L_X2Y125_SLICE_X0Y125_CO6),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D = CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_AMUX = CLBLL_L_X2Y116_SLICE_X1Y116_AO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_AMUX = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_BMUX = CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_CMUX = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_DMUX = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_AMUX = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_BMUX = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_AMUX = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_BMUX = CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_AMUX = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_BMUX = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_AMUX = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_AMUX = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_AMUX = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_CMUX = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_AMUX = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_BMUX = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_AMUX = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_AMUX = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_AMUX = CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B = CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C = CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D = CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_AMUX = CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D = CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B = CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D = CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B = CLBLL_L_X2Y128_SLICE_X1Y128_BO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C = CLBLL_L_X2Y128_SLICE_X1Y128_CO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D = CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_AMUX = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_AMUX = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_AMUX = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_AMUX = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_AMUX = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_BMUX = CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_AMUX = CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_CMUX = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_AMUX = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_AMUX = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_DMUX = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_AMUX = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_BMUX = CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_AMUX = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_CMUX = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_AMUX = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_AMUX = CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_AMUX = CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_AMUX = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_AMUX = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_AMUX = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_BMUX = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_AMUX = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_AMUX = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_AMUX = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_BMUX = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_AMUX = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A2 = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A3 = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A4 = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A5 = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B1 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B2 = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B3 = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B4 = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B5 = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B6 = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C1 = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C2 = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C4 = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C5 = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C6 = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = 1'b1;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A1 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B1 = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B3 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B5 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B6 = CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C2 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C5 = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C6 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D2 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D3 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D4 = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D6 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A2 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A5 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B2 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C1 = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C2 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D1 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D2 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D4 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D6 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A1 = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A4 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B2 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C2 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C3 = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C5 = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C6 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A2 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A3 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A4 = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A5 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A6 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B1 = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B2 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B3 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B5 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B6 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C1 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C5 = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C6 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D1 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D2 = CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D3 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D4 = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D6 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A6 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A2 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A3 = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A4 = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A5 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A6 = CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C6 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D6 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A2 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A4 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C2 = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C3 = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C4 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C6 = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D1 = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B1 = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B2 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B4 = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B5 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B6 = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C3 = CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C4 = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C5 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C2 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D2 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D3 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D6 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A1 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A2 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A3 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A4 = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A6 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B1 = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B3 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B4 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B5 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B6 = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D3 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D4 = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D5 = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B6 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C1 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C3 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A4 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B1 = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B5 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C1 = CLBLL_L_X2Y116_SLICE_X1Y116_AO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C2 = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C3 = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C4 = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C6 = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D1 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D2 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D3 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D4 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D6 = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A4 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B4 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C1 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C2 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C5 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C6 = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A2 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A5 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B5 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B6 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C3 = CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_D = LIOB33_X0Y121_IOB_X0Y121_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A1 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A3 = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A4 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B2 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B3 = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B4 = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A2 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A4 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B1 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B2 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B3 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B4 = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C1 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C2 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C3 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C5 = CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C6 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D2 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D3 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D6 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B1 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B2 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B3 = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B4 = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B6 = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C1 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D3 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D4 = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D5 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A2 = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A3 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A4 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A5 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A6 = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B2 = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B3 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B4 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B5 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B6 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C4 = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C5 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C6 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D2 = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D3 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D4 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D5 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D6 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A1 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A2 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A3 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A4 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A5 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A6 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B2 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B3 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B4 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B5 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B6 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C1 = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C2 = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C3 = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C4 = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C5 = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C6 = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D2 = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D3 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D4 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D5 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D6 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A1 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A4 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A6 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B1 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B5 = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B6 = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C6 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A6 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B2 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B4 = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B5 = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B6 = CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C1 = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C4 = CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C5 = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C6 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A5 = CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
endmodule
