module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CLK;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AMUX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BMUX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AQ;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BMUX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CLK;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_AMUX;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_BO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_BO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_CO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_DO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_AO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_BO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_BO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_CLK;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_CO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_DO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AMUX;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BMUX;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CMUX;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AMUX;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_AMUX;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_BO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_BO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_CO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_CO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_DO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_DO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_AO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_AO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_BO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_BO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_CLK;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_CO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_CO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_DO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_CO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_DO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_AO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_BO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_CO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_DO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_AMUX;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_BO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_CO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_DO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_AMUX;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_BO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_BO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_CO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_CO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_DO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_BO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_DO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AMUX;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_BO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_CO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_DO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A5Q;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CLK;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B5Q;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CLK;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C5Q;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CLK;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CLK;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CLK;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C5Q;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CLK;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CLK;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CLK;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DMUX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CLK;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A5Q;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CLK;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CLK;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CLK;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B5Q;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CLK;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B5Q;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BMUX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CLK;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CLK;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CLK;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AMUX;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CMUX;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5Q;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5Q;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B5Q;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B5Q;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AMUX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C5Q;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CMUX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A5Q;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B5Q;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D5Q;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AMUX;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D5Q;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DMUX;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A5Q;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AMUX;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AMUX;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BMUX;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CLK;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CLK;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CLK;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CMUX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CLK;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AMUX;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CLK;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_DO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AMUX;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AX;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BMUX;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CE;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CLK;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CMUX;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_SR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CLK;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CLK;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D5Q;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DMUX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CLK;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A5Q;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AMUX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CLK;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DMUX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CLK;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CLK;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DMUX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CLK;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DMUX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CLK;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AMUX;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CMUX;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_DO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CLK;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CMUX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_DO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CLK;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CMUX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DMUX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CE;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CLK;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_SR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CLK;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AMUX;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A5Q;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C5Q;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CE;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_SR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B5Q;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BMUX;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B5Q;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BMUX;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CE;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_SR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AMUX;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AMUX;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AMUX;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_AO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_AO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_BO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_BO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_CO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_CO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_DO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_DO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_AO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_BO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_BO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_CO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_CO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_DO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_DO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AMUX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CMUX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B5Q;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CLK;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CLK;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A5Q;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AMUX;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AX;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A5Q;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CLK;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D5Q;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CLK;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BMUX;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A5Q;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CLK;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CLK;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DMUX;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CLK;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CLK;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CE;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CLK;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_SR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CLK;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CLK;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_DO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CLK;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_DO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_BO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CLK;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_DO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_AO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_AO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_BO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_BO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_DO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_DO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CLK;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_DO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_BO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_DO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_DO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CLK;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CLK;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_DO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AMUX;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AX;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BMUX;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CE;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CLK;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_SR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AMUX;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CMUX;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AMUX;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CLK;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_DO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CLK;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CMUX;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_DO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CLK;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_DO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AQ;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CLK;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_CO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_DO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_AO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_AO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_BO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_BO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_CO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_CO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_DO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_DO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_AO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_AO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_BO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_BO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_CO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_CO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_DO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_DO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CLK;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CLK;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CLK;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DMUX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BMUX;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CLK;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CMUX;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AMUX;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_AMUX;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_AO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_BO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_BO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_CO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_CO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_DO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AMUX;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_BO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_DO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_DO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AMUX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CMUX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CLK;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CLK;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A5Q;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CLK;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CLK;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CLK;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CLK;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C5Q;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CMUX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D5Q;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A5Q;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666600cc00cc)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_ALUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_BO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbbfffbfffb)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbbfffffff3)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff3ffffffbb)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLL_L_X2Y126_SLICE_X1Y126_DO6),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0545004400440044)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_ALUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X1Y122_CO5),
.Q(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.Q(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.Q(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000500000c0d0c0c)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_DLUT (
.I0(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I1(LIOB33_X0Y63_IOB_X0Y63_I),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_DQ),
.I5(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88000000c8c0c0c0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_AQ),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc000c0ff600060)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_BLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X2Y123_SLICE_X1Y123_AQ),
.I5(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0cc00cc0fcc00)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_AQ),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I5(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff01ff01ff01ff55)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y123_SLICE_X0Y123_BO5),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.I4(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I5(CLBLL_L_X2Y123_SLICE_X0Y123_BO6),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ffffffaaaaffff)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbffffeffffff)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_ALUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.Q(CLBLL_L_X2Y123_SLICE_X1Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff3fff0)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y123_SLICE_X0Y123_AO5),
.I2(CLBLL_L_X2Y124_SLICE_X1Y124_CO6),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_AQ),
.I5(CLBLL_L_X2Y122_SLICE_X1Y122_DO6),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff000050dc)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_CLUT (
.I0(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I2(LIOB33_X0Y67_IOB_X0Y68_I),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_AO6),
.I4(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_BO6),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f50000fffdfffd)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff50ff5050505050)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_ALUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccccccdd)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_DLUT (
.I0(CLBLL_L_X2Y125_SLICE_X0Y125_DO6),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.I2(1'b1),
.I3(CLBLL_L_X2Y128_SLICE_X0Y128_CO6),
.I4(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.I5(CLBLM_R_X3Y124_SLICE_X3Y124_CO6),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_DO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000a003b000a)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_CLUT (
.I0(LIOB33_X0Y69_IOB_X0Y70_I),
.I1(CLBLL_L_X2Y123_SLICE_X0Y123_BO6),
.I2(CLBLL_L_X2Y125_SLICE_X0Y125_BO6),
.I3(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_CO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000000)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(LIOB33_X0Y67_IOB_X0Y68_I),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_BO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffaff7fff7ff)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_AO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y124_SLICE_X1Y124_AO6),
.Q(CLBLL_L_X2Y124_SLICE_X1Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffafafafe)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_DLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_BO6),
.I1(CLBLL_L_X2Y126_SLICE_X1Y126_CO6),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_DO6),
.I3(CLBLL_L_X2Y128_SLICE_X0Y128_CO6),
.I4(CLBLL_L_X2Y125_SLICE_X0Y125_BO5),
.I5(CLBLL_L_X2Y127_SLICE_X1Y127_DO6),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_DO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00330000003b000a)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_CLUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_AQ),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I4(LIOB33_X0Y57_IOB_X0Y58_I),
.I5(CLBLL_L_X2Y123_SLICE_X0Y123_BO6),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_CO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f020f00000202)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_BLUT (
.I0(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I1(CLBLL_L_X2Y123_SLICE_X0Y123_BO6),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I3(CLBLL_L_X2Y124_SLICE_X0Y124_AO5),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(LIOB33_X0Y57_IOB_X0Y57_I),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_BO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heccccccc20000000)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_ALUT (
.I0(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_AQ),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.I4(CLBLL_L_X2Y126_SLICE_X1Y126_AQ),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_AO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffffffbfffff)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X2Y125_SLICE_X0Y125_CO6),
.I4(CLBLL_L_X2Y124_SLICE_X0Y124_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00585058000a0a0a)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbbff08000800)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffffff08020800)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffccee)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_DLUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_DO6),
.I2(1'b1),
.I3(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I4(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.I5(CLBLL_L_X2Y124_SLICE_X1Y124_BO6),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000200)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_CLUT (
.I0(CLBLL_L_X2Y124_SLICE_X0Y124_AO6),
.I1(CLBLL_L_X2Y125_SLICE_X0Y125_CO6),
.I2(CLBLL_L_X2Y125_SLICE_X0Y125_BO5),
.I3(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.I5(CLBLL_L_X2Y126_SLICE_X0Y126_AO5),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_BLUT (
.I0(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.I1(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I2(CLBLL_L_X2Y125_SLICE_X0Y125_CO6),
.I3(CLBLL_L_X2Y126_SLICE_X0Y126_AO5),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_DO6),
.I5(CLBLL_L_X2Y123_SLICE_X0Y123_CO6),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffffffffbff)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0203020302000200)
  ) CLBLL_L_X2Y126_SLICE_X0Y126_DLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.I1(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I2(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.O5(CLBLL_L_X2Y126_SLICE_X0Y126_DO5),
.O6(CLBLL_L_X2Y126_SLICE_X0Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000000)
  ) CLBLL_L_X2Y126_SLICE_X0Y126_CLUT (
.I0(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_CO6),
.I3(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I4(CLBLL_L_X2Y124_SLICE_X0Y124_AO6),
.I5(CLBLL_L_X2Y125_SLICE_X0Y125_CO6),
.O5(CLBLL_L_X2Y126_SLICE_X0Y126_CO5),
.O6(CLBLL_L_X2Y126_SLICE_X0Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffbff)
  ) CLBLL_L_X2Y126_SLICE_X0Y126_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_AO6),
.I2(CLBLL_L_X2Y125_SLICE_X0Y125_CO6),
.I3(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I4(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.I5(CLBLL_L_X2Y126_SLICE_X0Y126_AO5),
.O5(CLBLL_L_X2Y126_SLICE_X0Y126_BO5),
.O6(CLBLL_L_X2Y126_SLICE_X0Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffff00080002)
  ) CLBLL_L_X2Y126_SLICE_X0Y126_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y126_SLICE_X0Y126_AO5),
.O6(CLBLL_L_X2Y126_SLICE_X0Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y126_SLICE_X1Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y126_SLICE_X1Y126_AO6),
.Q(CLBLL_L_X2Y126_SLICE_X1Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdfcfdfc)
  ) CLBLL_L_X2Y126_SLICE_X1Y126_DLUT (
.I0(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.I1(CLBLL_L_X2Y128_SLICE_X1Y128_CO6),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_BO6),
.I3(CLBLL_L_X2Y126_SLICE_X1Y126_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y126_SLICE_X5Y126_BO6),
.O5(CLBLL_L_X2Y126_SLICE_X1Y126_DO5),
.O6(CLBLL_L_X2Y126_SLICE_X1Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000000000000)
  ) CLBLL_L_X2Y126_SLICE_X1Y126_CLUT (
.I0(CLBLL_L_X2Y125_SLICE_X0Y125_CO6),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_CO6),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.I3(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I4(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I5(CLBLL_L_X2Y124_SLICE_X0Y124_AO6),
.O5(CLBLL_L_X2Y126_SLICE_X1Y126_CO5),
.O6(CLBLL_L_X2Y126_SLICE_X1Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7fffffff3)
  ) CLBLL_L_X2Y126_SLICE_X1Y126_BLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_CO6),
.I1(CLBLL_L_X2Y126_SLICE_X0Y126_BO6),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_BO6),
.I3(CLBLL_L_X2Y128_SLICE_X1Y128_BO6),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_CO6),
.O5(CLBLL_L_X2Y126_SLICE_X1Y126_BO5),
.O6(CLBLL_L_X2Y126_SLICE_X1Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff505050505050)
  ) CLBLL_L_X2Y126_SLICE_X1Y126_ALUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y126_SLICE_X1Y126_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_DQ),
.O5(CLBLL_L_X2Y126_SLICE_X1Y126_AO5),
.O6(CLBLL_L_X2Y126_SLICE_X1Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff2)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_DLUT (
.I0(CLBLL_L_X2Y126_SLICE_X1Y126_AQ),
.I1(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I2(CLBLL_L_X2Y126_SLICE_X0Y126_DO6),
.I3(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I4(CLBLL_L_X2Y128_SLICE_X0Y128_DO6),
.I5(CLBLL_L_X2Y127_SLICE_X0Y127_BO6),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_DO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888cccc88f8ccfc)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y61_I),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_CO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(LIOB33_X0Y55_IOB_X0Y55_I),
.I5(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_BO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202020202ff0202)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(CLBLL_L_X2Y125_SLICE_X0Y125_BO6),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I3(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I4(LIOB33_X0Y59_IOB_X0Y59_I),
.I5(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_AO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff4fffffff4f4)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_DLUT (
.I0(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I2(CLBLM_R_X3Y128_SLICE_X2Y128_AO5),
.I3(CLBLL_L_X2Y123_SLICE_X0Y123_AO6),
.I4(CLBLM_R_X3Y123_SLICE_X3Y123_DO6),
.I5(LIOB33_X0Y65_IOB_X0Y66_I),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_DO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdfffffffc)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_CLUT (
.I0(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.I1(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.I2(CLBLL_L_X2Y128_SLICE_X1Y128_DO6),
.I3(CLBLL_L_X2Y124_SLICE_X0Y124_CO6),
.I4(CLBLL_L_X2Y127_SLICE_X0Y127_AO6),
.I5(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_CO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_BO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_ALUT (
.I0(CLBLL_L_X2Y128_SLICE_X1Y128_DO6),
.I1(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.I2(CLBLL_L_X2Y127_SLICE_X0Y127_AO6),
.I3(CLBLL_L_X2Y127_SLICE_X1Y127_BO6),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_CO6),
.I5(CLBLL_L_X2Y124_SLICE_X0Y124_CO6),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_AO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000102200001000)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_DLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLL_L_X2Y125_SLICE_X0Y125_BO6),
.I5(LIOB33_X0Y71_IOB_X0Y71_I),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_DO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002000)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLL_L_X2Y125_SLICE_X0Y125_BO6),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_CO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000c0c5d0c)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_BLUT (
.I0(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I1(LIOB33_X0Y67_IOB_X0Y67_I),
.I2(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_BO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbffffbffff)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200020002020000)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I2(CLBLL_L_X2Y129_SLICE_X1Y129_AO5),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_DO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff4f4fff4)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_CLUT (
.I0(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.I2(CLBLM_R_X3Y128_SLICE_X2Y128_DO6),
.I3(LIOB33_X0Y67_IOB_X0Y67_I),
.I4(CLBLL_L_X2Y123_SLICE_X0Y123_AO6),
.I5(CLBLM_R_X3Y129_SLICE_X2Y129_BO6),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_CO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeefffffffe)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_BLUT (
.I0(CLBLM_R_X3Y128_SLICE_X2Y128_DO6),
.I1(CLBLL_L_X2Y128_SLICE_X0Y128_BO6),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_BO6),
.I4(CLBLM_R_X3Y128_SLICE_X2Y128_BO6),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_BO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffffffbfffff)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_ALUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_DO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_CO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_BO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_AO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_DO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_CO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_BO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffddff33ff33)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_AO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfc69966996)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_AO5),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_AO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_BO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2aaa2a200ff0000)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.I2(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_A5Q),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaefaa00004500)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.I5(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f000f101f000)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_BLUT (
.I0(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000cacacaca)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_ALUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_AO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffffefafffff)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_DLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbbbbbbbc0000000)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DQ),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac0c0aaaa30c0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y122_SLICE_X5Y122_AO5),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaffaa0faa0f)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I2(LIOB33_X0Y53_IOB_X0Y53_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_CO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heecceecceac0eac0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0eef0eef0ee)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_CLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_CQ),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I5(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ddfff0f08800)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5550ccccfff0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_ALUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_C5Q),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.I3(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X5Y122_BO5),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X5Y122_AO6),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffffffffffffff)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_DLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_DQ),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1333200033330000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_CLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_CO6),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_B5Q),
.I5(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c5c5fffff000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_BLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.I1(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff1212125f5f5f5f)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_CO6),
.I2(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X4Y123_CO5),
.Q(CLBLL_L_X4Y123_SLICE_X4Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X4Y123_AO6),
.Q(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X4Y123_BO6),
.Q(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X4Y123_CO6),
.Q(CLBLL_L_X4Y123_SLICE_X4Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000a0c0a0c)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_DQ),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaccaacc)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_CLUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faaffaa0caacc)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I1(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefcfefcaa00aa00)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.I2(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_D5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_AO6),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_CO6),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044554400)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_DLUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I5(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f3f4f007030400)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_CQ),
.I5(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3333aaaa0000)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_BLUT (
.I0(CLBLL_L_X4Y123_SLICE_X5Y123_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff80ff0000800000)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_ALUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_B5Q),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_D5Q),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.Q(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.Q(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_DLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_CO6),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_CO5),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffffccdfdfdf)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000000f000f)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_D5Q),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_C5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000800000008)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_ALUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_C5Q),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_CO5),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_AO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_BO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_CO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hceffceffcececece)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_CO6),
.I2(CLBLL_L_X2Y125_SLICE_X0Y125_AO6),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888fa50fa50)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0003300cc)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000320032)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d5d5d5d0c0c0c0c)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_DLUT (
.I0(CLBLL_L_X2Y125_SLICE_X0Y125_AO6),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_CQ),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff77ff55ff33ff00)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_CLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_CO5),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.I2(1'b1),
.I3(CLBLL_L_X4Y123_SLICE_X4Y123_DO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_BLUT (
.I0(CLBLL_L_X2Y125_SLICE_X1Y125_DO6),
.I1(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_DO6),
.I3(CLBLL_L_X2Y125_SLICE_X1Y125_BO6),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_CO6),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3f3aaaac0c0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_ALUT (
.I0(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_A5Q),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X5Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff4f4fff4)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_DLUT (
.I0(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_DO6),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_BO6),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fdf55dd0fcf00cc)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_CLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_CO5),
.I1(CLBLL_L_X4Y122_SLICE_X5Y122_B5Q),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I3(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I5(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000080000)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_D5Q),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfa0c0afcfa0c0a)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55550000f5f5f0f0)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_DLUT (
.I0(CLBLL_L_X2Y125_SLICE_X0Y125_AO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_DO5),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f555f550f000f00)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_CLUT (
.I0(CLBLL_L_X2Y125_SLICE_X0Y125_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y122_SLICE_X7Y122_DQ),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h73735050ff73ff50)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_CO6),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I4(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22f222f2ffff22f2)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_ALUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.I5(CLBLM_R_X3Y125_SLICE_X2Y125_CO6),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X5Y126_AO6),
.Q(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff4fff44)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_DLUT (
.I0(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.I3(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.I4(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_CO6),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f550f00dfddcfcc)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I5(CLBLL_L_X2Y125_SLICE_X0Y125_AO6),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00aaaaa0a0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_ALUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_B5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_AO5),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_AO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_BO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffffffffff7)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfffffffeff)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haacfaaffaac0aa00)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_BLUT (
.I0(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00f0f0aaaa)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_CQ),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.I3(RIOB33_X105Y127_IOB_X1Y127_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_AO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0eef000f0ee)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_BLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_B5Q),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfe0032fefe3232)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_ALUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I3(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I5(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_BO6),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff44fffffff4)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_DLUT (
.I0(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_CO6),
.I4(CLBLL_L_X4Y129_SLICE_X4Y129_DO6),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_DO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000000)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_CO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa0caa0faa0c)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_BO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8dddd8888888)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I4(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_AO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_BO5),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_AO6),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_BO6),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030ffff30303030)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_CQ),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_DO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffee)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_CLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_A5Q),
.I5(CLBLL_L_X4Y129_SLICE_X5Y129_BO6),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_CO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f40404cfc0cfc0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_BO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4455445544504450)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_ALUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_CQ),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_AO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_BO5),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_AO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_CO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_DLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0055554444)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ccaaccaa)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_BLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3cccaaaacccc)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_ALUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.I3(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y130_SLICE_X3Y130_CQ),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_AO6),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdd)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_B5Q),
.I2(1'b1),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_CO6),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_CQ),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_CLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_B5Q),
.I3(CLBLL_L_X4Y129_SLICE_X4Y129_B5Q),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_A5Q),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_BLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_CQ),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_B5Q),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I3(CLBLM_L_X8Y128_SLICE_X10Y128_B5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_B5Q),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0cccc)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_AO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_BO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_CO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_DO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff28ff2828282828)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_DLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_DO6),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_DO5),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f8f8f822888888)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_DO6),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_A5Q),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I5(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6fcf0f066cc0000)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_BLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_AO6),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_DO6),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf0fcc00fcf0cc00)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_DO6),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_AO6),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_CO6),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffa)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_DLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I3(CLBLL_L_X4Y124_SLICE_X5Y124_CQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_A5Q),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0707ffff7777ffff)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_CLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.I5(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_BLUT (
.I0(CLBLM_R_X3Y126_SLICE_X2Y126_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_B5Q),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_DO6),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_DO6),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_A5Q),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I5(CLBLL_L_X4Y130_SLICE_X4Y130_CQ),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_AO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8cc000000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ce0202020202)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0e2c0c0e2c0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_CO6),
.I4(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fe32cc00dc10)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_AO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_BO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_CO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_DO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00ff00f0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000ee00ee)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fe04fe04)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_BQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc5055550000)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_CO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h010104010b0b0e0b)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_DLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_A5Q),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfff50a00)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc55cc00cc55)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_DO6),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b88888b8b8)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_BO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050005)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffffffbffff)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_DO6),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f000f0cc)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_C5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc0acc00)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ff66ffff66ff66)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff77bbddee)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_CLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_A5Q),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003f00ff002e00)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_BLUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_DO6),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I5(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccffcc00)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_CO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_DO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaa1100baaa1000)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y123_SLICE_X14Y123_A5Q),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88dd88888888)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff504000005040)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0ffaaaa0000)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_ALUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I3(CLBLM_L_X8Y123_SLICE_X11Y123_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_BO6),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008400840000)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_DO6),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_CO6),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_DQ),
.I5(CLBLM_L_X8Y123_SLICE_X11Y123_BO6),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fdf000000000ff)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X2Y126_SLICE_X1Y126_DO6),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000fcfc)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_CQ),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafefe00005454)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_BO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff00ffffe0e0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_DQ),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd88888fff00000)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0006060c0c)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0055555050)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_ALUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_D5Q),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_C5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha353a353a303a353)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_BLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_DQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_CO6),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_DO6),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303f303f000f000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_CO5),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_BO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_CO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa880000aacc0000)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_AO5),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf000ff00aaaa)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_C5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01ab01ba10ba10)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_AO5),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a0a0ffcc0000)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I2(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_BO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c33c3cc30000)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_DQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc00c8c8c8c8)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff540054ff540054)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc4ffc8c4c4c8c8)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_ALUT (
.I0(CLBLM_L_X8Y126_SLICE_X11Y126_CO6),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hab81aaa0aaa0aaa0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaeaaa20004)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000003300330)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcfcfc00)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I4(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbf000005050000)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_DLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_CO5),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000320022)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_CLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_CO5),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcd0101cece0202)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_BLUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5550cccc5550)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_ALUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.Q(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.R(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_DLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfecffcc13203300)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_CLUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_AO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc88cc88cc88dc18)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05050505afafafaf)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_ALUT (
.I0(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_AO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_BO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfcfdfccdcccdcc)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_CO6),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h669999995aa5a5a5)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_BQ),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_DO6),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_AO6),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_DO6),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888b8b8b8b8888)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_CO6),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff323200003232)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_ALUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_CQ),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_BO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_CO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_DO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c0c5c5c0c5c0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafcf80f0a0c08)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afc0cfc0c)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_BLUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_A5Q),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd888d888d8)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_D5Q),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_BO5),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_BO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303030303030)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8dddddd8d888888)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_DO6),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeae0404dd88dd88)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I4(CLBLM_R_X11Y128_SLICE_X15Y128_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fa50aa00fa50)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_BO5),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_CO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_DLUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f2f1f404020104)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y129_SLICE_X14Y129_CQ),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_DO6),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaf0f0ccf0cc)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_BLUT (
.I0(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_A5Q),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc0fcc00cc00)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33c3cc3c33c)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffdd0000fddd)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_CO5),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I2(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_D5Q),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fa50ee44ea40)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_CO6),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff60ff6000600060)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_ALUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_DO6),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_DQ),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_CO5),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_AO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_BO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_CO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c333f0f0a0a0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_DLUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccaaccaacc)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_CLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I1(RIOB33_X105Y125_IOB_X1Y126_I),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0003030c0c)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccfa05050505)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeeffffffff)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_DLUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I1(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdffffffff)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_CLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000010)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_CQ),
.I1(CLBLM_R_X11Y129_SLICE_X14Y129_CQ),
.I2(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I3(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I4(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000004000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_ALUT (
.I0(CLBLM_L_X8Y129_SLICE_X11Y129_DO6),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_BO6),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_CO6),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_BO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_CO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_DO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaefeae04045404)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5e4f5a0a0e4a0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_B5Q),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff50d8000050d8)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_BLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf50055005500)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_BO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000800000003)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee44440f0f0000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hce02cd01ce02cd01)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5500ccccf5a0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_ALUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_DQ),
.I2(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_CO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0a0a005050000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_DLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33003300)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0afafafa0ac)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_BLUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88b888b8bbbb8888)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_ALUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I5(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555f5555ffff)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.I1(1'b1),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555fffffff7)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_CLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c000a000a0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_BLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccf0ccaaccaa)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I5(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_AO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb055bb552f662277)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_BLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I3(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0000f05a)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_ALUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_DO6),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I2(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I3(CLBLM_L_X8Y132_SLICE_X10Y132_BO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.R(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333000033333333)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_DO6),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000f5f5f5f5)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y135_SLICE_X16Y135_AO5),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h020e010d020e010d)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_A5Q),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f3c0f3f3)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff50ff5000500050)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_A5Q),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000e000ff1fff0ff)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000054155550541)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_CLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_AO6),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f3c0f3f3)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdf0020dddddddd)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_ALUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4f0b4f0f0f0f0f0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_DLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c287d7d28)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_CLUT (
.I0(CLBLM_R_X3Y126_SLICE_X2Y126_CO6),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_A5Q),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.I5(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeefffffe01ff00)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_BLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300f0d2f0f0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_ALUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb04fb04ff00ff00)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_DLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000efff10ffff)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_A5Q),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fe5403030303)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd02ff0022222222)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccd8cccc)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_AO6),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I5(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe02fd0102fe01fd)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I2(CLBLM_R_X3Y126_SLICE_X2Y126_CO6),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_BO5),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_D5Q),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_DO6),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.I5(CLBLM_L_X10Y120_SLICE_X13Y120_CO6),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa47748bb8)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_ALUT (
.I0(CLBLM_R_X11Y122_SLICE_X15Y122_A5Q),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_AO6),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_DQ),
.I5(CLBLM_R_X3Y126_SLICE_X2Y126_CO6),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_BO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_CO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc333c333c)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000aa00aa)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_CLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_A5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0fff0cc)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdecdec00120120)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_ALUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I5(CLBLM_L_X10Y127_SLICE_X13Y127_C5Q),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_BO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f06030603)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_DLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_CO5),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_AO5),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc9cccc0f0fffff)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff45ff4500450045)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_BLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_DO6),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fb0400003333)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_CO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_DO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fffa5550)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_DQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fefe5454)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_B5Q),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacff0ff000)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_BLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafffcaaaa0030)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_ALUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00550055cc883377)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_DLUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_DO6),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y126_SLICE_X1Y126_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffccf0f0aa88)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0a0a0aca0a0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_CO6),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0c0c0c0c0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_DQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_B5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_CLUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_D5Q),
.I1(CLBLM_L_X8Y123_SLICE_X11Y123_DO6),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_DO6),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_CQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_DO6),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_CQ),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff03ff3000030030)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_CO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0f202f202)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_DLUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4e48888dd88)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_DQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcac0c00055ffff)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_BLUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_A5Q),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32dc10fe32dc10)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_ALUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_CO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_DO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccedccde00210012)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_A5Q),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_B5Q),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecececc02020200)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c0c0ff00c0c0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00fc30)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_ALUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccccf0a0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0e0e00000e0e)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000eee0eee0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_BLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaafff0ffc0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_CO6),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffaa)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_DLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I5(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc0000f0f0aaaa)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_CLUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0cfcfc0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_DQ),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_CO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefecc32323200)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300330033)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_D5Q),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fbfb00000b0b)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_CLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_DO6),
.I5(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808f808cfcfc0c0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafff0ccc0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_B5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I3(CLBLM_L_X12Y125_SLICE_X17Y125_DQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_AO5),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_BO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000fffe)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_DLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_DO6),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_CO6),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_BQ),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_CLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I1(CLBLM_L_X10Y127_SLICE_X13Y127_C5Q),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I5(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afacafacafac)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I5(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fa50e4e4e4e4)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X13Y126_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.Q(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa88aa888aa8aa88)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_AO6),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_C5Q),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555655fffff3f3)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_CLUT (
.I0(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccff0000cc0000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_DQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfccccc30300000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_BO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_BO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_CO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050505090505)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_DLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcfcac0c0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0e4e4a0a0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_DQ),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ec20aaaaa0a0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_D5Q),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_CO5),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_AO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_BO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_CO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_DO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f033f011f011)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_DLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_CO6),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacaa0afa0a0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_CLUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_C5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d8d8d8d88888888)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddcdddc11101110)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_ALUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_CO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_AO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_AO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00001010f3f3f3f3)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_DLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_BO6),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(1'b1),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff500050ffddffdd)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y129_SLICE_X15Y129_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0ffdd)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_R_X11Y130_SLICE_X15Y130_BO6),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaafffff0c0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_ALUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_DO5),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_BO6),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_DO6),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0fafa0a0a)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_DLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_A5Q),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11cc00dd11cc00)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0d1d1c0c0e2e2)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_BLUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y128_SLICE_X13Y128_CQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_CQ),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2c0aaaaaa00)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_AO5),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_BO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_DO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00a000a0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_DQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c0c5c5c0c5c0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_AO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaba1010baba1010)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3a0a0fa0afa0a)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_ALUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_A5Q),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I4(CLBLM_R_X11Y129_SLICE_X15Y129_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_DO5),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_AO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_BO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0aaaacccc)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_DLUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I2(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fe0ef000fe0e)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_CLUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00ff00cc)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_BLUT (
.I0(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454feaa5400)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_CO6),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_CO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_AO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_BO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_CO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc3333c333)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLM_L_X10Y130_SLICE_X13Y130_DO6),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fff0ff00555055)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_DO6),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff15ff1400150014)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I2(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_DO6),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_A5Q),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8dddddddddddd)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I2(CLBLM_R_X11Y130_SLICE_X15Y130_BO6),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.Q(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0088110008881000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_DLUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00001040efbf)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33001300cc00ec00)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_AO6),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30333033f0ff3033)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.I5(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_CO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3ccc3ccc33cc33)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555dddd05050d0d)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.I5(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f9f009f0f0f000f)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_BLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_BO6),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I5(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd00ddddd0000dddd)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.I5(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ffffffd5ffffff)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_DLUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f500f500ff00f7)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_DO6),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ef00cf00ef00ef)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_AO5),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4303400003030000)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f03030f0f0303)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb00bbbbb0000bbbb)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_CO6),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.I5(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_AO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_CO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_DO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa5555aaaa5595)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_DLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_CO6),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_DO6),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_BO5),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_DO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h333333333c333333)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_DO6),
.I3(CLBLM_L_X12Y122_SLICE_X16Y122_CO6),
.I4(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_CO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010001000500050)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_BLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I3(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_BO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cca0000000f0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.I1(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_AO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_DO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_BO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_AO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X16Y121_BO6),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h333f333f333f333f)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_BO6),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_DQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0000ff55)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_CLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_L_X12Y122_SLICE_X17Y122_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f000f101f000)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_DQ),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_CO6),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefcfbf3aa00aa00)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_ALUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_DQ),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_BO6),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X16Y122_AO6),
.Q(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X16Y122_BO6),
.Q(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y125_SLICE_X17Y125_CQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0b00000044)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_BO6),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcc0c0000cc0c)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0ffcc00a000cc)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X17Y122_AO6),
.Q(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.Q(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X17Y122_CO6),
.Q(CLBLM_L_X12Y122_SLICE_X17Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haac0aaffaac0aa00)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_CLUT (
.I0(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I1(CLBLM_L_X12Y122_SLICE_X17Y122_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I5(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eeaaf0f0aaaa)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_CO6),
.I1(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaffaaf0aaf0)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff3f3fcfc)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_DO6),
.I3(1'b1),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I5(CLBLM_R_X11Y123_SLICE_X15Y123_DO6),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_DO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ff66ffff66ff66)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_CLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I1(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y125_SLICE_X17Y125_BQ),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_CO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd5da808fd5da808)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_BLUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_BO5),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_BO6),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_BO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc8cc800000000)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_DO6),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_BO5),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_DO6),
.I5(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_AO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X17Y123_AO6),
.Q(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffefffe)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_DLUT (
.I0(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I1(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I3(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_DO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa55555511)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_DO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_AO5),
.I4(CLBLM_L_X12Y123_SLICE_X17Y123_DO6),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_CO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333233)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_BLUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_DO6),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I2(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_DO6),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I5(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_BO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8ffffffaa)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_ALUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I3(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_AO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_DQ),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.R(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6fff6fffff6fff6)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_DLUT (
.I0(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_CO6),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000300010303030)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_CLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080088000000)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_BLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff0004040404)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_A5Q),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X17Y124_AO6),
.Q(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X17Y124_BO6),
.Q(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X17Y124_CO6),
.Q(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X17Y124_DO6),
.Q(CLBLM_L_X12Y124_SLICE_X17Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafc00)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_DLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I2(CLBLM_L_X12Y124_SLICE_X17Y124_DQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd800d8ff500050)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I1(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.I2(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf0fafa0c000a0a)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_BLUT (
.I0(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.I1(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddd8888888d8)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.I2(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_L_X12Y124_SLICE_X17Y124_DQ),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_DO5),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_DO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccaaaaff00)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_DLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_B5Q),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I3(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_DO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f6f00600)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_CLUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_CO5),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_CO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfbccbbf0f00000)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_BLUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_BO5),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I3(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_CO6),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_BO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fcaaaa0000)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_ALUT (
.I0(CLBLM_L_X12Y125_SLICE_X17Y125_DQ),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_BO6),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_AO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X17Y125_AO6),
.Q(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X17Y125_BO6),
.Q(CLBLM_L_X12Y125_SLICE_X17Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X17Y125_CO6),
.Q(CLBLM_L_X12Y125_SLICE_X17Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X17Y125_DO6),
.Q(CLBLM_L_X12Y125_SLICE_X17Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafeaa00005400)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_DQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_DO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacf0faaaac000)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_CLUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_CQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_CO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00fef40e04)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_DQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_BO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aafcaaf0aafc)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_AO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_DO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_BO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8bbbbb800ff0000)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_DLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_A5Q),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0caaffaa0caa00)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_CLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_CQ),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.I5(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff55f0f0ff44)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_CQ),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cddc0110)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_ALUT (
.I0(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_DO5),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_AO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafabfafeafabfafe)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_DLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I2(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I3(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haeffaeaa04550400)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ee22ee22)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdcde0000dcde)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_ALUT (
.I0(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I3(CLBLM_L_X12Y128_SLICE_X17Y128_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_AO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_BO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_CO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010001000000010)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_DLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_A5Q),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888bb88bb8b)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_CLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I4(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I5(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0c0caaaaff00)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_BLUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_CQ),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0330aaaa0030)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_ALUT (
.I0(CLBLM_L_X12Y124_SLICE_X17Y124_DQ),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I3(CLBLM_L_X12Y124_SLICE_X16Y124_AO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X17Y127_AO6),
.Q(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X17Y127_BO6),
.Q(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X17Y127_CO6),
.Q(CLBLM_L_X12Y127_SLICE_X17Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000200)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_DLUT (
.I0(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I2(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I4(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaccaaf0aaf0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_CQ),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505fd0df000f808)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_CQ),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff454100004541)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X13Y126_SLICE_X19Y126_CO6),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_AO6),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_BO6),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_CO6),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_DO6),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0f00fc00)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_DLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_DO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa03030c03)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_CLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_CO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ff55eb41)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.I2(CLBLM_R_X13Y128_SLICE_X19Y128_BO6),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_BO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfcccfc00300030)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y128_SLICE_X17Y128_CO6),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_AO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0810081008108800)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_DLUT (
.I0(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I2(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I4(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I5(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_DO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeafbebebebebebe)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_CLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I3(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.I4(CLBLM_L_X12Y128_SLICE_X17Y128_DO6),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_CO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555551554555)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_BLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_DO5),
.I3(CLBLM_R_X13Y126_SLICE_X18Y126_CQ),
.I4(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I5(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_BO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005533333f7f)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_ALUT (
.I0(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_CO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X16Y129_AO6),
.Q(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.Q(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hce003b000a00ce00)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_DLUT (
.I0(CLBLM_L_X12Y129_SLICE_X16Y129_CO5),
.I1(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_DO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h020000000a0a0000)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_CLUT (
.I0(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I1(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_CO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfccccc33320000)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_BLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I4(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_BO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555eafa4050)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I5(CLBLM_L_X12Y129_SLICE_X16Y129_CO6),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_AO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X17Y129_AO6),
.Q(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.Q(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0a7757eeee0000)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_DLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I4(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_DO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001aa01cbca41ca)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_CLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I2(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f099cc)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_BLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_DO6),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I2(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_BO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb88b888bb888b)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.I5(CLBLM_L_X12Y128_SLICE_X17Y128_BO6),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_AO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.R(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.Q(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000050)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_DLUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000010000)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_CLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffffff)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I5(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccffccf0ccf0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fdd11cc00)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffcfffffefef)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.Q(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaffc0ffeaeac0c0)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_CLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I2(LIOB33_X0Y51_IOB_X0Y51_I),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0e0a0c000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_BLUT (
.I0(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.I4(LIOB33_X0Y53_IOB_X0Y53_I),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00f3f3ffff)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.Q(CLBLM_R_X3Y122_SLICE_X2Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55a0c0c0c0c)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_CLUT (
.I0(CLBLL_L_X2Y126_SLICE_X1Y126_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55c3c93c36)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd1ff0000d10000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_ALUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_CO6),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.Q(CLBLM_R_X3Y122_SLICE_X3Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff77ff77ffffffff)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_DLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_AQ),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1100000015000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_BLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hed21cc00fc30cc00)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_ALUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I5(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff05ff01ffffffff)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_DLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_C5Q),
.I1(CLBLL_L_X2Y124_SLICE_X1Y124_AQ),
.I2(LIOB33_X0Y53_IOB_X0Y53_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_CLUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000a000c)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_BLUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X2Y123_SLICE_X0Y123_BO5),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeefffe)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_ALUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_CO6),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_BO6),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_BO6),
.I4(CLBLL_L_X2Y125_SLICE_X0Y125_AO6),
.I5(CLBLM_R_X3Y123_SLICE_X2Y123_CO6),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1011100000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_DLUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I1(CLBLL_L_X2Y123_SLICE_X0Y123_BO5),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccce000affff000a)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I3(CLBLL_L_X2Y125_SLICE_X0Y125_BO6),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_CQ),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500454405000500)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_BLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.I2(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_ALUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h888faaaf8888aaaa)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_DLUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_C5Q),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_AO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff2fffffff22)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_CLUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I1(CLBLL_L_X2Y125_SLICE_X0Y125_AO6),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.I3(CLBLL_L_X2Y124_SLICE_X0Y124_BO6),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_DO6),
.I5(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1100110011005150)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_BLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I2(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_ALUT (
.I0(CLBLM_R_X3Y123_SLICE_X3Y123_DO6),
.I1(CLBLM_R_X3Y123_SLICE_X2Y123_BO6),
.I2(CLBLM_R_X3Y126_SLICE_X2Y126_AO6),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.I4(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_DO6),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3fff0fff33ff00)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.I2(CLBLM_R_X3Y125_SLICE_X2Y125_CO6),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_DO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff50ffffff5050)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_CLUT (
.I0(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.I4(CLBLM_R_X3Y125_SLICE_X3Y125_BO6),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aacceef0fafcfe)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_BLUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.I4(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I5(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000101033003310)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I2(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I5(CLBLL_L_X2Y125_SLICE_X0Y125_BO6),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y125_SLICE_X2Y125_AO6),
.Q(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd00df0fdd00dd00)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_DLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_BO5),
.I5(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbffffdfff)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f7ffffffffefef)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(1'b1),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfcccfc00f000f0)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.I3(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fcfcfafafefe)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_DLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_CLUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_DO6),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_DO6),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_DO6),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_CO6),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_BO6),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h03000b0a03000300)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I4(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffffffffeff)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecececeffceffce)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_DLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.I1(CLBLM_R_X3Y128_SLICE_X3Y128_CO6),
.I2(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000100)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_CLUT (
.I0(CLBLL_L_X2Y126_SLICE_X1Y126_BO6),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I4(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I5(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300030057550300)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_BLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I1(CLBLL_L_X2Y125_SLICE_X0Y125_BO6),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.I5(CLBLM_R_X3Y129_SLICE_X2Y129_AO6),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff10551010)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_ALUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I2(LIOB33_X0Y65_IOB_X0Y66_I),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_BO5),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I5(CLBLM_R_X3Y128_SLICE_X2Y128_AO5),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff50ffffff50ff50)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_DLUT (
.I0(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.I1(1'b1),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_CO6),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_CO6),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000330050507350)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_CLUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_BO5),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.I4(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I5(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_BLUT (
.I0(CLBLL_L_X2Y127_SLICE_X0Y127_DO6),
.I1(CLBLL_L_X4Y126_SLICE_X4Y126_AO6),
.I2(CLBLL_L_X2Y125_SLICE_X1Y125_BO6),
.I3(CLBLL_L_X4Y126_SLICE_X4Y126_CO6),
.I4(CLBLL_L_X4Y128_SLICE_X4Y128_DO6),
.I5(CLBLM_R_X3Y125_SLICE_X3Y125_DO6),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbffffffbfff)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfefffffcfe)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_DLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I1(CLBLM_R_X3Y128_SLICE_X2Y128_CO6),
.I2(CLBLM_R_X3Y126_SLICE_X2Y126_BO6),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_CO6),
.I4(CLBLM_R_X3Y128_SLICE_X3Y128_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_DO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_CLUT (
.I0(CLBLM_R_X3Y129_SLICE_X2Y129_CO6),
.I1(CLBLL_L_X2Y125_SLICE_X1Y125_BO6),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_DO6),
.I4(CLBLL_L_X2Y127_SLICE_X1Y127_CO6),
.I5(CLBLM_R_X3Y126_SLICE_X2Y126_DO6),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_CO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cae0caeffff0cae)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_DQ),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_CO6),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_CO6),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_BO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_ALUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.I1(CLBLL_L_X2Y125_SLICE_X1Y125_BO6),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_DO6),
.I3(CLBLL_L_X2Y127_SLICE_X1Y127_AO6),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_AO6),
.I5(CLBLL_L_X2Y126_SLICE_X0Y126_CO6),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_AO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafafaffaafffa)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_DLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_AO6),
.I1(1'b1),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_CO6),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_DO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff22fffffff2)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_CLUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_CO6),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_CO6),
.I4(CLBLM_R_X3Y128_SLICE_X3Y128_DO6),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_CO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefffefe)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_BLUT (
.I0(CLBLM_R_X3Y127_SLICE_X3Y127_DO6),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_DO6),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_DO6),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_DO6),
.I4(CLBLL_L_X2Y125_SLICE_X1Y125_CO6),
.I5(CLBLM_R_X3Y127_SLICE_X3Y127_CO6),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_BO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30ba30baffff30ba)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_CO6),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I5(CLBLM_R_X3Y125_SLICE_X2Y125_CO6),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_AO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011000100100000)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_DLUT (
.I0(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_DO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000a000accce)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I5(CLBLM_R_X3Y129_SLICE_X2Y129_AO6),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_CO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000c05050000)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_BLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I2(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I4(CLBLM_R_X7Y127_SLICE_X9Y127_DQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_BO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfdfdf500f500)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_AO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'habffaaff03030000)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(LIOB33_X0Y65_IOB_X0Y65_I),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_DO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000cc005000dc)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_CLUT (
.I0(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_CQ),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_CO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d888888888888)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_DO5),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(CLBLM_R_X3Y128_SLICE_X3Y128_AO5),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_BO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffafffaf0a000a00)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(1'b1),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_AO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200000002505)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_DLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLM_R_X3Y128_SLICE_X3Y128_AO5),
.I4(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I5(CLBLL_L_X2Y129_SLICE_X1Y129_AO6),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400040007030400)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_CLUT (
.I0(CLBLM_R_X3Y129_SLICE_X2Y129_AO5),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.I5(CLBLL_L_X2Y129_SLICE_X1Y129_AO6),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0d5c0ccccddcc)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_BLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_C5Q),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_AO6),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfffdffff3fff3)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X3Y129_AO6),
.Q(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X3Y129_BO6),
.Q(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeeffffffff)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(1'b1),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_CQ),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f5f5e4e4a0a0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_CQ),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888bb88888)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X2Y130_AO6),
.Q(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fff00000f0f0)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X3Y130_DO6),
.Q(CLBLM_R_X3Y130_SLICE_X3Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.Q(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.Q(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X3Y130_CO6),
.Q(CLBLM_R_X3Y130_SLICE_X3Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaac0c00000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_DLUT (
.I0(RIOB33_X105Y127_IOB_X1Y127_I),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f606f000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_CLUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaaeeaa3c00cc00)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_BLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_CQ),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_CQ),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdecceecc5a00aa00)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_ALUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_CQ),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_AO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_BO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_DLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_CLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa003000c0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_BLUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000480048)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I3(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_CO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000fdfd)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_DLUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cacacacac)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_CLUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0aaf0ccf088)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f044cccc0000)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff030f33ff030f)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.I2(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.I3(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I4(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff20ff0020200000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.I5(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h030f0f0fa3afafaf)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_DO6),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X2Y126_SLICE_X1Y126_DO6),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_CO6),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88eeee2222)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_BO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_CO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f8f8f8f8f8f8f8f)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_DLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000fc00)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_CLUT (
.I0(CLBLL_L_X2Y124_SLICE_X1Y124_AQ),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_CQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaa0caaccaa0c)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_BLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_B5Q),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff84ff8400840084)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_ALUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_AO5),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_BO6),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc44cc00cc)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I5(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0fff8fffcff)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_CLUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I5(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafa0050aaea0040)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_A5Q),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44fff0004400f0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_BO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_CO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50ee44ee44)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_DQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0eeeeee00)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_BLUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_DO6),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeceeecaaa0aaa0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_ALUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_BO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_CO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_DO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa30fc3030)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_DLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32ee22ce02ee22)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.I3(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I5(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaafcaa00aa0c)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_BLUT (
.I0(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_CO6),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfefe00003232)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_ALUT (
.I0(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I5(CLBLL_L_X4Y123_SLICE_X4Y123_CQ),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_BO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_CO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_DO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05500550)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y124_SLICE_X5Y124_C5Q),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_DO6),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000e0e0e0e)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_CLUT (
.I0(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I3(1'b1),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0ccf0aaf0cc)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbff5155eaaa4000)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I5(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_AO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_BO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_CO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000000)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f0fc0003000c)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_BQ),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdd0011ddcc1100)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_D5Q),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_DO6),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd800d8ffd800d8)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_ALUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_BO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_CO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_DO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaf0aaf0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaafaa05000500)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00f0f0cccc)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0aaccccf0aa)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdfdfdfccdfdfdf)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_DLUT (
.I0(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.I3(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.I4(CLBLL_L_X2Y126_SLICE_X1Y126_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a00000aaaa0000)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_CLUT (
.I0(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_DO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_BLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_DO6),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I3(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc55cc00cc50)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_CO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000032023202)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05ff55ae04ee44)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.I5(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefef4f40e0e0404)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3f3aaaac0c0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_ALUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_DLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h32223000ffffffff)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_CLUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_CO5),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aabfbfbf)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I4(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I5(CLBLM_R_X5Y125_SLICE_X7Y125_CO6),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff007777ff007070)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_CO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafc00)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_DLUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I1(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_DQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffee00ee00ee00)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_CLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_DQ),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fcfc0f000c0c)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I5(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfaaafaaa)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_ALUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_BO6),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_DO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_BO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5e400330033)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_A5Q),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff005500ee0044)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfe0ef000f000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y122_SLICE_X7Y122_DQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fa000afcfa0c0a)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_CO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_DO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd8dd8dddd8)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff88ff88ff888888)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0fffaaaa0ccc)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0c00aaaa0c00)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_ALUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff22fff2ff22fff2)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_DLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_DO5),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_CO6),
.I4(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808080000080000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_DO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303f303f303f000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeeeeee50444444)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_BQ),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_AO5),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_DO5),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_CO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_DO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f00ff00aaaa)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_DLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00cb00cb00cb)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_CLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000acacacac)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_DQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I3(1'b1),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cfcfc0c0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_ALUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_CO5),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_CO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffffffffffff)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_DLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0aaffaa00)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_CLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X2Y126_SLICE_X1Y126_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf00c00fcfc0c0c)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_C5Q),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccfff000cc00f0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_DO5),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_BO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_CO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_DO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f03300aaaaf0f0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_DLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500feae5404)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff000c0c)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaaff00)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_ALUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_CQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_BO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeeeeeeeeeee)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0a00000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_CLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_D5Q),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcff0c0ffcf00c00)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I5(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00fafa0a0a)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_ALUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaffaaffaa)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_DLUT (
.I0(CLBLL_L_X4Y129_SLICE_X4Y129_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0e0e00000e0e)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_CLUT (
.I0(CLBLL_L_X4Y129_SLICE_X4Y129_B5Q),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ffcc3300)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_BLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I4(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haeea0cc0aeea0cc0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_DO6),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_BO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccfcffcecfcec)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_DLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haabfbfbfc0000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_CLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_CQ),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f606fc0c)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_BLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_AO6),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cfcfc0c0c0c5)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a000a000a000)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_DLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0b1a0e4a0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_DO6),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaaf888faaaf888)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0aa000000aa0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_ALUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_CO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500eeee4444)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0c0c0cfc0c0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffc0f0c0f0c)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_B5Q),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_BO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111111100000000)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fe00ff01010000)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_CLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc5cfcacfc5cfca)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_BLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_DO6),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacac5cac0c0c0c0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_ALUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_AO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaafaaaa)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_CLUT (
.I0(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I5(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccdcffffff00)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_BLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_CO6),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I3(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.I4(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00fcfc)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X9Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cac0cac0cac0c0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_CO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_CO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000003)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.I2(CLBLL_L_X2Y126_SLICE_X1Y126_DO6),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaafe00540054)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fcfc0c0c)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_A5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000033303330)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_CO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_BO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f700f500f700f5)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0e455445544)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000a0aff000808)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccfc00330030)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000ebaa4100)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_CO6),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.I5(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00000ee00)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_B5Q),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffa0afc0cf808)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc50ccf0ccfaccf0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0f3f0f000f00)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbfffa)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffb300)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccdcccc00010000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(CLBLM_R_X5Y126_SLICE_X7Y126_CQ),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4040404000000000)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa030caaaa0c0c)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_CLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_D5Q),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0eef000f044)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeecaaa0eeecaaa0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_ALUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_CO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a05000000a05)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_DLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_D5Q),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_DO6),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000ff0fc5c5c0c0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_C5Q),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_D5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f606f000f606)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_CO6),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fc000000fc)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_BO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_CO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_DO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fe54fe54fe54)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_DQ),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11aa00bb11aa00)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f404f404)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeecaaa0eeecaaa0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_ALUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_DLUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_DO5),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00a000ff00c0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_CLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaacc00ff0fff)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_BLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c8c8c8cccccc00)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_B5Q),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_CO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_DLUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafaaa50005000)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f606f606)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cfc0c0cf)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8888dddd8888d)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.I3(CLBLM_L_X10Y126_SLICE_X13Y126_CO5),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0ffac00ff0000)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_AO6),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0cfcfc0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_AO5),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f5fa050a)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffffffffffffff)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I4(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4e4a0a0e4e4)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fcfc0f000c0c)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5050ccccff50)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dbe7dbe7dbe7dbe)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_DLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_DQ),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_A5Q),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000008000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_CLUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_DQ),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_DQ),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_DO6),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_DO6),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f303f000fc0c)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ccccfafa)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_A5Q),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_DQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_DO5),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaff00ccccf0f0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_DLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d8f0d8f0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_CLUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I3(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aafcaafcaafc)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_BLUT (
.I0(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I5(CLBLM_L_X12Y122_SLICE_X16Y122_BQ),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacaca0afafafa0af)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_ALUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_BO5),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaff55005500)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_DQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f0000c0c0caca)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22fccc3000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I4(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa30aa33aa30)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_ALUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_B5Q),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_BO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_CO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_DO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0aaaa00cc)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f033cc)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y129_SLICE_X10Y129_DO5),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01ab01ba10ba10)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0aaf0ccf0aa)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_ALUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_CO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_DO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00fafafa)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_DLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_DQ),
.I3(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f044444444)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I2(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb888888bb8888)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0f3f3c0c0f3c0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_BO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880000000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_A5Q),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_CLUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_A5Q),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_DO6),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.I5(CLBLM_R_X7Y128_SLICE_X8Y128_DO6),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcaca0000caca)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_BLUT (
.I0(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff003030)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y128_SLICE_X8Y128_CO6),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_CO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdfff)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_DLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff08ff0800080008)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c5c0c0c5c5c0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_BO5),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fc30cc00fc30)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_BO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44000000baba1010)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h54550000fcff0000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c0c0ff00c0c0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_D5Q),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd888dd88d888d888)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_CO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_BO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h005500ff00fc00fc)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_DLUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef00e000f000f00)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_CLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_D5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafcf0fafafcf0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_BLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.I2(CLBLM_L_X8Y129_SLICE_X11Y129_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaafff0ffc0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_ALUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_A5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BO6),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaaabaaa10001000)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_DQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff5aa0a0a0a0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_A5Q),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f606fc0c)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_BLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_CQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_DQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_AO6),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f077fff0f0ffff)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_CO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_DO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888d8d8d8d8)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dddd8888)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y144_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a0a3a0ff0ff000)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_BLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_BQ),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc00ccf5cca0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_ALUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I1(CLBLL_L_X2Y126_SLICE_X1Y126_AQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_BO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffaaaa)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_DLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaafaa05000500)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c0c0c5c5c0c0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_BLUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff44e4000044e4)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_ALUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5522ddaf507788)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_DLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555f5555555755)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_DO6),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_DO6),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafc0a0cfaff0a0f)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_DO6),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.I4(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05555f0f00000)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_ALUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.I1(1'b1),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h08a208a28888888a)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_DO6),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fc000001fc00000)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I4(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_DO6),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddcccdc11100010)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_DO6),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00fe44444545)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_DO6),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003030ff003030)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff77ffc0c00000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y139_IOB_X1Y140_I),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.I4(RIOB33_X105Y141_IOB_X1Y141_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c000000aaaaaaa6)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_ALUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_AO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000000404040)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f000f044f000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_DQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00eeaaeca0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_ALUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_AO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_BO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_DLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.I5(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h050503030505030c)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_CLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afa0afaf)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_BLUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_DQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdf0020eeffeeff)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_BO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f00000f0f0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd5ff55aad5aa55)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_CLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h666666666c666666)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_BLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I3(CLBLM_L_X12Y122_SLICE_X16Y122_CO6),
.I4(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_DO6),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5ad25a5a)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_DO6),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_CO6),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I4(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_DO6),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeeee0e0e0e0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_DO6),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0311030003220333)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_CLUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_BO6),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_CQ),
.I2(CLBLM_L_X10Y128_SLICE_X13Y128_DQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff002222f0f0ff55)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_BLUT (
.I0(RIOB33_X105Y119_IOB_X1Y119_I),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aa30aaf0aa30)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_ALUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_B5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X15Y121_AO6),
.Q(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X15Y121_BO6),
.Q(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaaaaabbaa)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_DQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c3f00002e1d)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_CLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_A5Q),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_DQ),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heac0eac0eac0ffc0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_BLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_BO6),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffc00fc00fc)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_BO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff3000ffff30)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_DO6),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300000f5a)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_CLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_BO6),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0e000eff0e000e)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_BLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafff0ccc0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_B5Q),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X15Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X15Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaaa55aa5555aa)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa55aa5a55aa55a)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_CLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y125_SLICE_X17Y125_BQ),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0906090606090609)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_BLUT (
.I0(CLBLM_R_X11Y122_SLICE_X15Y122_DO6),
.I1(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y122_SLICE_X15Y122_CO6),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe3232ccfe0032)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.I4(CLBLM_R_X11Y128_SLICE_X15Y128_DQ),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_DO5),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_AO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_BO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccaaffaa00)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_DLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaffaa00)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0003030c0c)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_DO6),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I4(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8ffcc3300)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_ALUT (
.I0(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I4(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X15Y123_AO6),
.Q(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X15Y123_BO6),
.Q(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X15Y123_CO6),
.Q(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ffff6666ffff66)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_DLUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I1(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff54ff5400540054)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000f0c0f0c)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I4(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d580d580)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_ALUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I3(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_CO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_DLUT (
.I0(CLBLM_R_X11Y123_SLICE_X15Y123_BQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafacafaca0a0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_CLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_CO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fc0cf000fc0c)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaafa00550050)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00f3000000f3)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff54ff5400540054)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000c0aac0aa)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_BLUT (
.I0(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I4(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc005acccc0000)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_ALUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_CO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_A5Q),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_CO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_DO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd8ffd8ffd8ff88)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_C5Q),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_DQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_DO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00af05af05aa00)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_BO5),
.I5(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0ef000eeee0000)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_B5Q),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00ccccfa50)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X15Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X15Y125_BO6),
.Q(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X15Y125_CO6),
.Q(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00aa00ff00aa)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafae0504aaaa0000)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_CO6),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000060c060c)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_BLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_DO6),
.I1(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffaaffccffa0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_ALUT (
.I0(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_D5Q),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_CO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_BQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb8888888888)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5a0f5a0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_B5Q),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22ee22fc30)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_CQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_AO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_BO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_CO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_DO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaeaaaaafaea)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f4f5f405040504)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000e0eff000000)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_BLUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_DQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff0033dcfe1032)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I3(CLBLM_L_X10Y126_SLICE_X13Y126_CO6),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_DO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffe0ff00ffe0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffee000000ee)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_CLUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaa00fcfc0000)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_BLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_CQ),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff5000550050)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_ALUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X15Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X15Y127_BO6),
.Q(CLBLM_R_X11Y127_SLICE_X15Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X15Y127_CO6),
.Q(CLBLM_R_X11Y127_SLICE_X15Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffcc0000fafa)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_CQ),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafc00)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_CLUT (
.I0(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_CQ),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_DO6),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404f404f404)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfd3131fefe3232)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_ALUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I5(CLBLM_L_X12Y127_SLICE_X16Y127_DO6),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_BO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_CO5),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_AO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_BO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffddffdc)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_DLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I1(CLBLM_R_X11Y129_SLICE_X14Y129_DO6),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.I3(CLBLM_L_X10Y130_SLICE_X13Y130_BO6),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccaaaa)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2c0aaaaaa00)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_CQ),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aafcaa00aafc)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_BO6),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_AO6),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_DO6),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454feaa5400)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_DO6),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_DQ),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_DQ),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c5c5caca)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I1(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X11Y128_SLICE_X15Y128_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf80a08aa88aa88)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_DQ),
.I4(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdff0000fdff)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLM_R_X11Y130_SLICE_X15Y130_BO6),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y128_SLICE_X12Y128_B5Q),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_AO6),
.Q(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_BO6),
.Q(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_CO6),
.Q(CLBLM_R_X11Y129_SLICE_X14Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffffffdffff)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_DLUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_DO6),
.I1(CLBLM_R_X11Y130_SLICE_X15Y130_CO6),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_DO6),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff055000000550)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y128_SLICE_X13Y128_AO5),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0f3f3)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_DO6),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe400e4ffe400e4)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_ALUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_CQ),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y129_SLICE_X15Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X15Y129_AO6),
.Q(CLBLM_R_X11Y129_SLICE_X15Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X15Y129_BO6),
.Q(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X15Y129_CO6),
.Q(CLBLM_R_X11Y129_SLICE_X15Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5544554455555050)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I1(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_DQ),
.I4(CLBLM_R_X11Y129_SLICE_X15Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f022222222)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_CLUT (
.I0(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32fe32fe32fe32)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000fc00)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_ALUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_CO6),
.I2(CLBLM_R_X11Y129_SLICE_X15Y129_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_AO6),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_BO6),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_CO6),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555577775555)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaac0f0c0c0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f30000f3f3)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.I5(CLBLM_L_X10Y130_SLICE_X13Y130_BO6),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff00fdfd)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLM_R_X11Y130_SLICE_X15Y130_BO6),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X15Y130_AO6),
.Q(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff5)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_DQ),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc50cc00cc50)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fff7fffffffff)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_DLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000effbffff)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.I2(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30003030ff00ffff)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_BO6),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80aac0ff08aa0cff)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500550055550000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_DLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_CO6),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_CO6),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_CLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000cf3ff0008f7)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_BLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_CO6),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_CO6),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333310033333333)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_DO6),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I5(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.Q(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.R(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f3c0f3c0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_AO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_BO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_CO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_DLUT (
.I0(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.I2(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.I3(CLBLM_L_X12Y122_SLICE_X17Y122_CQ),
.I4(CLBLM_L_X12Y125_SLICE_X17Y125_CQ),
.I5(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_DO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff008f8fff008080)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y125_SLICE_X17Y125_CQ),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_CO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd8ff5000d80050)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb3ff8000b30080)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_DQ),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_AO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X19Y123_AO6),
.Q(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X19Y123_BO6),
.Q(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X19Y123_CO6),
.Q(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_DO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f5a0a0a0f5a0)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y123_SLICE_X19Y123_CQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_CO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffd5800000d580)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I1(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_BO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf30b03f8f00800)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_ALUT (
.I0(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_CQ),
.I5(CLBLM_L_X12Y122_SLICE_X17Y122_CQ),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_AO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y124_SLICE_X18Y124_AO6),
.Q(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_DO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_CO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_BO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a0a0ff00cccc)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.I2(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_AO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_DO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_CO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_BO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_AO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y125_SLICE_X18Y125_AO6),
.Q(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fffa0f0a)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_ALUT (
.I0(CLBLM_R_X13Y128_SLICE_X18Y128_AO6),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_AO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_DO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_CO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_BO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_AO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.Q(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X18Y126_BO6),
.Q(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X18Y126_CO6),
.Q(CLBLM_R_X13Y126_SLICE_X18Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.Q(CLBLM_R_X13Y126_SLICE_X18Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5500ccccf5a0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_DLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_DQ),
.I3(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05500f0f0dd88)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_CLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_CQ),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_CO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcefe0232cece0202)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_BO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0eff0e000e000e)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_AO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X19Y126_AO6),
.Q(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_DO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffffffff)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_CLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_CQ),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_CO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_BLUT (
.I0(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.I5(CLBLM_R_X13Y129_SLICE_X19Y129_CO6),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_BO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfa5150fbfa5150)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I2(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_AO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.Q(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.R(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000100)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_DLUT (
.I0(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6633666366666666)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_CLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_DO6),
.I3(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_DQ),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f7ffff55000000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_BLUT (
.I0(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_AO5),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h222222330f0f0f0e)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_ALUT (
.I0(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_AO5),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I4(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ffffffffffffff)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_DLUT (
.I0(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I1(CLBLM_R_X13Y129_SLICE_X19Y129_CO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000100)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_CLUT (
.I0(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h333399cc33339ccc)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_BLUT (
.I0(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_AQ),
.I2(CLBLM_R_X13Y126_SLICE_X19Y126_BO6),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_CQ),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I5(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5151404051514040)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_ALUT (
.I0(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_AQ),
.I2(CLBLM_R_X13Y126_SLICE_X19Y126_BO6),
.I3(1'b1),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_DLUT (
.I0(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_DO5),
.I5(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_DO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_CLUT (
.I0(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_DO5),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_CO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f4f0f0f0f4fc)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_BLUT (
.I0(CLBLM_R_X13Y128_SLICE_X18Y128_DO6),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.I2(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I4(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_CO6),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_BO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc23dc33cc03fc)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_ALUT (
.I0(CLBLM_R_X13Y128_SLICE_X18Y128_DO6),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_CQ),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I4(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_CO6),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_AO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.Q(CLBLM_R_X13Y128_SLICE_X19Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333fffb3333ffff)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_DLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I5(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_DO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002200000020)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_CLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I1(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I5(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_CO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5151555151555555)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_BLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.I2(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I4(CLBLM_R_X13Y129_SLICE_X19Y129_CO6),
.I5(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_BO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888ddd88888ddd8)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_BO6),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_AO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.Q(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.Q(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fe2222fff22222)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_DLUT (
.I0(CLBLM_R_X13Y129_SLICE_X18Y129_CO5),
.I1(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I3(CLBLM_R_X13Y129_SLICE_X18Y129_CO6),
.I4(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_A5Q),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_DO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habab11bb000000f0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_CLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_CO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0aaf000f0aa)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_BLUT (
.I0(CLBLM_R_X13Y129_SLICE_X18Y129_DO6),
.I1(1'b1),
.I2(CLBLM_R_X13Y128_SLICE_X19Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_CO6),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_BO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ef45fe54)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_BO6),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_AO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y129_SLICE_X19Y129_AO6),
.Q(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff11ff33ff51ff)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_DLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I3(CLBLM_R_X11Y129_SLICE_X15Y129_CQ),
.I4(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_DO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h444c000000000000)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_CLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I4(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_CO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666665665666)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_BLUT (
.I0(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_DO5),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I5(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_BO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afacafac)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_ALUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y129_SLICE_X19Y129_BO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_AO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.Q(CLBLM_R_X13Y132_SLICE_X18Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_DO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_CO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_BO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0fff0f0)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_DO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_CO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_AO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y122_SLICE_X56Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y122_SLICE_X56Y122_DO5),
.O6(CLBLM_R_X37Y122_SLICE_X56Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y122_SLICE_X56Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y122_SLICE_X56Y122_CO5),
.O6(CLBLM_R_X37Y122_SLICE_X56Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y122_SLICE_X56Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y122_SLICE_X56Y122_BO5),
.O6(CLBLM_R_X37Y122_SLICE_X56Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f0000)
  ) CLBLM_R_X37Y122_SLICE_X56Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.I3(1'b1),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X37Y122_SLICE_X56Y122_AO5),
.O6(CLBLM_R_X37Y122_SLICE_X56Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y122_SLICE_X57Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y122_SLICE_X57Y122_DO5),
.O6(CLBLM_R_X37Y122_SLICE_X57Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y122_SLICE_X57Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y122_SLICE_X57Y122_CO5),
.O6(CLBLM_R_X37Y122_SLICE_X57Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y122_SLICE_X57Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y122_SLICE_X57Y122_BO5),
.O6(CLBLM_R_X37Y122_SLICE_X57Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y122_SLICE_X57Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y122_SLICE_X57Y122_AO5),
.O6(CLBLM_R_X37Y122_SLICE_X57Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_ALUT (
.I0(RIOB33_X105Y139_IOB_X1Y139_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafffff0f0f)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0fff0fff0f)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I4(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfffff0f0ffff)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_DO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_CO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_BO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_AO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_DO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_CO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_BO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeeffeeffee)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_ALUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(1'b1),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_AO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfffff0f0ffff)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y123_SLICE_X1Y123_BO5),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_R_X11Y123_SLICE_X14Y123_D5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X11Y123_SLICE_X14Y123_DQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X10Y123_SLICE_X13Y123_DQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X8Y129_SLICE_X10Y129_C5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X3Y130_SLICE_X3Y130_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X7Y126_SLICE_X8Y126_D5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X11Y128_SLICE_X14Y128_C5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X2Y124_SLICE_X1Y124_AQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X3Y130_SLICE_X3Y130_CQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X3Y130_SLICE_X3Y130_BQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y138_SLICE_X163Y138_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_R_X7Y137_SLICE_X8Y137_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_BO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLM_R_X37Y122_SLICE_X56Y122_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_R_X11Y125_SLICE_X15Y125_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_R_X11Y129_SLICE_X15Y129_DO6),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_R_X11Y129_SLICE_X15Y129_DO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_R_X11Y127_SLICE_X15Y127_DO6),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_R_X11Y127_SLICE_X15Y127_DO5),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_L_X8Y134_SLICE_X11Y134_AO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO6),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_R_X11Y125_SLICE_X15Y125_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_R_X11Y129_SLICE_X15Y129_DO6),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_R_X11Y129_SLICE_X15Y129_DO5),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_R_X11Y127_SLICE_X15Y127_DO6),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_R_X11Y127_SLICE_X15Y127_DO5),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X13Y132_SLICE_X18Y132_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X103Y176_SLICE_X163Y176_AO6),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X103Y176_SLICE_X163Y176_AO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X13Y132_SLICE_X18Y132_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_AMUX = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_AMUX = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_BMUX = CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_CMUX = CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_AMUX = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_CMUX = CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_DMUX = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_AMUX = CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_BMUX = CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B = CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C = CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_BMUX = CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B = CLBLL_L_X2Y124_SLICE_X0Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_AMUX = CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B = CLBLL_L_X2Y124_SLICE_X1Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D = CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_AMUX = CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_BMUX = CLBLL_L_X2Y125_SLICE_X0Y125_BO5;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_CMUX = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D = CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_AMUX = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B = CLBLL_L_X2Y126_SLICE_X0Y126_BO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C = CLBLL_L_X2Y126_SLICE_X0Y126_CO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D = CLBLL_L_X2Y126_SLICE_X0Y126_DO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_AMUX = CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A = CLBLL_L_X2Y126_SLICE_X1Y126_AO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B = CLBLL_L_X2Y126_SLICE_X1Y126_BO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C = CLBLL_L_X2Y126_SLICE_X1Y126_CO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B = CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D = CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A = CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B = CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C = CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D = CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B = CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D = CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_AMUX = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B = CLBLL_L_X2Y128_SLICE_X1Y128_BO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C = CLBLL_L_X2Y128_SLICE_X1Y128_CO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D = CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_AMUX = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B = CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D = CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A = CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B = CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C = CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D = CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_AMUX = CLBLL_L_X2Y129_SLICE_X1Y129_AO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_AMUX = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A = CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_AMUX = CLBLL_L_X4Y121_SLICE_X4Y121_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_DMUX = CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A = CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_CMUX = CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_DMUX = CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A = CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_AMUX = CLBLL_L_X4Y122_SLICE_X5Y122_AO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_BMUX = CLBLL_L_X4Y122_SLICE_X5Y122_B5Q;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_CMUX = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A = CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B = CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C = CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_CMUX = CLBLL_L_X4Y123_SLICE_X4Y123_C5Q;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C = CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_CMUX = CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_DMUX = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A = CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B = CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C = CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_CMUX = CLBLL_L_X4Y124_SLICE_X5Y124_C5Q;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A = CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C = CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_DMUX = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A = CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_DMUX = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A = CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B = CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_AMUX = CLBLL_L_X4Y127_SLICE_X4Y127_A5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_CMUX = CLBLL_L_X4Y127_SLICE_X4Y127_CO5;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_DMUX = CLBLL_L_X4Y127_SLICE_X4Y127_DO5;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A = CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B = CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C = CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D = CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_DMUX = CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A = CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B = CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D = CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_BMUX = CLBLL_L_X4Y128_SLICE_X5Y128_B5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_DMUX = CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A = CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_BMUX = CLBLL_L_X4Y129_SLICE_X4Y129_B5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A = CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C = CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A = CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B = CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_DMUX = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_AMUX = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_BMUX = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_CMUX = CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B = CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C = CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A = CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B = CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C = CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A = CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_AMUX = CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C = CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_DMUX = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A = CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_AMUX = CLBLM_L_X8Y121_SLICE_X11Y121_A5Q;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_DMUX = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A = CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C = CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D = CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A = CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B = CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_AMUX = CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_CMUX = CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A = CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_CMUX = CLBLM_L_X8Y123_SLICE_X10Y123_CO5;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A = CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_CMUX = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A = CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B = CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C = CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_AMUX = CLBLM_L_X8Y124_SLICE_X10Y124_AO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_CMUX = CLBLM_L_X8Y124_SLICE_X10Y124_C5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A = CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_CMUX = CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A = CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B = CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A = CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B = CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_AMUX = CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_BMUX = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CMUX = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A = CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B = CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A = CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B = CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C = CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D = CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A = CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B = CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_BMUX = CLBLM_L_X8Y127_SLICE_X11Y127_B5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A = CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B = CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C = CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D = CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_BMUX = CLBLM_L_X8Y128_SLICE_X10Y128_B5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A = CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B = CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C = CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A = CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C = CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D = CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_AMUX = CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_CMUX = CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_DMUX = CLBLM_L_X8Y129_SLICE_X10Y129_DO5;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A = CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B = CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C = CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D = CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A = CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C = CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_AMUX = CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_CMUX = CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_DMUX = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_DMUX = CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A = CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_AMUX = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_BMUX = CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A = CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_BMUX = CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A = CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B = CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A = CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B = CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_AMUX = CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A = CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A = CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_AMUX = CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_DMUX = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_AMUX = CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_BMUX = CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_AMUX = CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_BMUX = CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_CMUX = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A = CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B = CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A = CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_AMUX = CLBLM_L_X10Y121_SLICE_X13Y121_AO5;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_CMUX = CLBLM_L_X10Y121_SLICE_X13Y121_CO5;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_BMUX = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A = CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_AMUX = CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_DMUX = CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_BMUX = CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_CMUX = CLBLM_L_X10Y123_SLICE_X13Y123_C5Q;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_DMUX = CLBLM_L_X10Y123_SLICE_X13Y123_D5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A = CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B = CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_AMUX = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A = CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CMUX = CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A = CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_BMUX = CLBLM_L_X10Y125_SLICE_X13Y125_B5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A = CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_AMUX = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_BMUX = CLBLM_L_X10Y126_SLICE_X12Y126_B5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A = CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_CMUX = CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A = CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B = CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C = CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_AMUX = CLBLM_L_X10Y127_SLICE_X12Y127_AO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A = CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B = CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D = CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_CMUX = CLBLM_L_X10Y127_SLICE_X13Y127_C5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C = CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_AMUX = CLBLM_L_X10Y128_SLICE_X12Y128_A5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_BMUX = CLBLM_L_X10Y128_SLICE_X12Y128_B5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_CMUX = CLBLM_L_X10Y128_SLICE_X12Y128_CO5;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_DMUX = CLBLM_L_X10Y128_SLICE_X12Y128_DO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B = CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_AMUX = CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_DMUX = CLBLM_L_X10Y128_SLICE_X13Y128_D5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B = CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D = CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_AMUX = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A = CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B = CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_DMUX = CLBLM_L_X10Y129_SLICE_X13Y129_D5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A = CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_AMUX = CLBLM_L_X10Y130_SLICE_X12Y130_A5Q;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_AMUX = CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B = CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A = CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B = CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C = CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D = CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_AMUX = CLBLM_L_X12Y120_SLICE_X16Y120_AO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_BMUX = CLBLM_L_X12Y120_SLICE_X16Y120_BO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A = CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A = CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B = CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C = CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A = CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B = CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_CMUX = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A = CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B = CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C = CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A = CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B = CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_AMUX = CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A = CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C = CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D = CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_AMUX = CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_BMUX = CLBLM_L_X12Y124_SLICE_X16Y124_BO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_CMUX = CLBLM_L_X12Y124_SLICE_X16Y124_CO5;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A = CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B = CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C = CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_DMUX = CLBLM_L_X12Y125_SLICE_X16Y125_D5Q;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A = CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B = CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C = CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D = CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_AMUX = CLBLM_L_X12Y126_SLICE_X16Y126_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_DMUX = CLBLM_L_X12Y126_SLICE_X16Y126_DO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A = CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A = CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B = CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C = CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D = CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_DMUX = CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A = CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_DMUX = CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A = CLBLM_L_X12Y128_SLICE_X16Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B = CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C = CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D = CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A = CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B = CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C = CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D = CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_AMUX = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_CMUX = CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A = CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_CMUX = CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A = CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D = CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_CMUX = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_DMUX = CLBLM_L_X12Y129_SLICE_X17Y129_DO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A = CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B = CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C = CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D = CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D = CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A = CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D = CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D = CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_AMUX = CLBLM_L_X12Y135_SLICE_X16Y135_AO5;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D = CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_AMUX = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_AMUX = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_BMUX = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_CMUX = CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_DMUX = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_BMUX = CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_CMUX = CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_AMUX = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A = CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_BMUX = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D = CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_AMUX = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_BMUX = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B = CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_BMUX = CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C = CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D = CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B = CLBLM_R_X3Y128_SLICE_X2Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C = CLBLM_R_X3Y128_SLICE_X2Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D = CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_AMUX = CLBLM_R_X3Y128_SLICE_X2Y128_AO5;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C = CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D = CLBLM_R_X3Y128_SLICE_X3Y128_DO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_AMUX = CLBLM_R_X3Y128_SLICE_X3Y128_AO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B = CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D = CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_AMUX = CLBLM_R_X3Y129_SLICE_X2Y129_AO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_CMUX = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A = CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B = CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A = CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C = CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D = CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C = CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D = CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_AMUX = CLBLM_R_X3Y130_SLICE_X3Y130_A5Q;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_DMUX = CLBLM_R_X3Y130_SLICE_X3Y130_DO5;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B = CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A = CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_CMUX = CLBLM_R_X3Y131_SLICE_X3Y131_CO5;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_AMUX = CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CMUX = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_AMUX = CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A = CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_DMUX = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A = CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B = CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A = CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B = CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B = CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C = CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A = CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B = CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C = CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A = CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B = CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D = CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A = CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_BMUX = CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_CMUX = CLBLM_R_X5Y124_SLICE_X7Y124_CO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A = CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B = CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A = CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_AMUX = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_AMUX = CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_DMUX = CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A = CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B = CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A = CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B = CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A = CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B = CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_AMUX = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_DMUX = CLBLM_R_X5Y128_SLICE_X6Y128_D5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A = CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B = CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C = CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_CMUX = CLBLM_R_X5Y128_SLICE_X7Y128_C5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A = CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_DMUX = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A = CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B = CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_BMUX = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CMUX = CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A = CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B = CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A = CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B = CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C = CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B = CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_CMUX = CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A = CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A = CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C = CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_BMUX = CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_AMUX = CLBLM_R_X7Y120_SLICE_X8Y120_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_AMUX = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CMUX = CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_DMUX = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A = CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_CMUX = CLBLM_R_X7Y122_SLICE_X9Y122_C5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A = CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B = CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C = CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_AMUX = CLBLM_R_X7Y123_SLICE_X9Y123_AO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_BMUX = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A = CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B = CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A = CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B = CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_CMUX = CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A = CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C = CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_DMUX = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_AMUX = CLBLM_R_X7Y126_SLICE_X9Y126_A5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_BMUX = CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CMUX = CLBLM_R_X7Y126_SLICE_X9Y126_CO5;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_DMUX = CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A = CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D = CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_DMUX = CLBLM_R_X7Y127_SLICE_X8Y127_D5Q;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A = CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B = CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C = CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D = CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_DMUX = CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A = CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C = CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A = CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B = CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_AMUX = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CMUX = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_DMUX = CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A = CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_AMUX = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_CMUX = CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_DMUX = CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A = CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B = CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_AMUX = CLBLM_R_X7Y130_SLICE_X8Y130_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CMUX = CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A = CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_BMUX = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CMUX = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A = CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A = CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_BMUX = CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B = CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C = CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_AMUX = CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A = CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B = CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_AMUX = CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_CMUX = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_AMUX = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A = CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B = CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C = CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_CMUX = CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_BMUX = CLBLM_R_X11Y121_SLICE_X14Y121_B5Q;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A = CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_AMUX = CLBLM_R_X11Y122_SLICE_X15Y122_A5Q;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_AMUX = CLBLM_R_X11Y123_SLICE_X14Y123_A5Q;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_DMUX = CLBLM_R_X11Y123_SLICE_X14Y123_D5Q;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B = CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A = CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B = CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C = CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A = CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A = CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C = CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_BMUX = CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A = CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B = CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C = CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C = CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D = CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A = CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B = CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A = CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D = CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_BMUX = CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A = CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_DMUX = CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A = CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B = CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_AMUX = CLBLM_R_X11Y128_SLICE_X14Y128_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_BMUX = CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_CMUX = CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A = CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_AMUX = CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_BMUX = CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A = CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B = CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C = CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B = CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_DMUX = CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A = CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B = CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C = CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A = CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C = CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D = CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A = CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B = CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D = CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A = CLBLM_R_X13Y123_SLICE_X18Y123_AO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B = CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C = CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D = CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A = CLBLM_R_X13Y123_SLICE_X19Y123_AO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B = CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C = CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D = CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A = CLBLM_R_X13Y124_SLICE_X18Y124_AO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B = CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C = CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D = CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A = CLBLM_R_X13Y124_SLICE_X19Y124_AO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B = CLBLM_R_X13Y124_SLICE_X19Y124_BO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C = CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D = CLBLM_R_X13Y124_SLICE_X19Y124_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A = CLBLM_R_X13Y125_SLICE_X18Y125_AO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C = CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D = CLBLM_R_X13Y125_SLICE_X18Y125_DO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A = CLBLM_R_X13Y125_SLICE_X19Y125_AO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C = CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D = CLBLM_R_X13Y125_SLICE_X19Y125_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B = CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C = CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A = CLBLM_R_X13Y126_SLICE_X19Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B = CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C = CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D = CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_AMUX = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_BMUX = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D = CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_AMUX = CLBLM_R_X13Y127_SLICE_X19Y127_AO5;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_CMUX = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A = CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B = CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_AMUX = CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B = CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C = CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D = CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_CMUX = CLBLM_R_X13Y129_SLICE_X18Y129_CO5;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A = CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B = CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C = CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D = CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B = CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D = CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A = CLBLM_R_X37Y122_SLICE_X56Y122_AO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B = CLBLM_R_X37Y122_SLICE_X56Y122_BO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C = CLBLM_R_X37Y122_SLICE_X56Y122_CO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D = CLBLM_R_X37Y122_SLICE_X56Y122_DO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A = CLBLM_R_X37Y122_SLICE_X57Y122_AO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B = CLBLM_R_X37Y122_SLICE_X57Y122_BO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C = CLBLM_R_X37Y122_SLICE_X57Y122_CO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D = CLBLM_R_X37Y122_SLICE_X57Y122_DO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A = CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B = CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C = CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D = CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B = CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C = CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D = CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_AMUX = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A = CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B = CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C = CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D = CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B = CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C = CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D = CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_AMUX = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A = CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B = CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C = CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D = CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B = CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C = CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D = CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_AMUX = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A = CLBLM_R_X103Y176_SLICE_X162Y176_AO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B = CLBLM_R_X103Y176_SLICE_X162Y176_BO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C = CLBLM_R_X103Y176_SLICE_X162Y176_CO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D = CLBLM_R_X103Y176_SLICE_X162Y176_DO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B = CLBLM_R_X103Y176_SLICE_X163Y176_BO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C = CLBLM_R_X103Y176_SLICE_X163Y176_CO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D = CLBLM_R_X103Y176_SLICE_X163Y176_DO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_R_X11Y123_SLICE_X14Y123_D5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X11Y123_SLICE_X14Y123_DQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X3Y130_SLICE_X3Y130_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X3Y130_SLICE_X3Y130_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X10Y123_SLICE_X13Y123_DQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X13Y132_SLICE_X18Y132_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLM_R_X37Y122_SLICE_X56Y122_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X13Y132_SLICE_X18Y132_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C1 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C4 = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C5 = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C6 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B1 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A1 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A4 = CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A5 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A6 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B2 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B4 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B5 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B6 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C1 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_AX = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C2 = CLBLM_L_X10Y129_SLICE_X13Y129_D5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C5 = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A1 = CLBLL_L_X4Y130_SLICE_X4Y130_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A3 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A4 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A6 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B2 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B3 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B6 = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C2 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C4 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C5 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D3 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLM_R_X37Y122_SLICE_X56Y122_AO6;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D5 = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X13Y132_SLICE_X18Y132_AQ;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B1 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B2 = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B5 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A1 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A2 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A4 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A5 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A6 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B1 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B2 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B4 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B5 = CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B6 = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C1 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C2 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C3 = CLBLL_L_X4Y130_SLICE_X4Y130_CQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D1 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D3 = CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D4 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A2 = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A3 = CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A4 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A5 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B1 = CLBLL_L_X4Y130_SLICE_X4Y130_CQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B3 = CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B4 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B5 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C1 = CLBLL_L_X4Y129_SLICE_X4Y129_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C2 = CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D1 = CLBLL_L_X4Y129_SLICE_X4Y129_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C3 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C5 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D2 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D3 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A2 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A4 = CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A6 = CLBLM_L_X8Y127_SLICE_X11Y127_B5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B2 = CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B4 = CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A3 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A4 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A5 = CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C2 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B1 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B2 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B4 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B5 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B6 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D2 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C1 = CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C2 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C3 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C4 = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C5 = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C6 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D4 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A1 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A2 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A3 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A4 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A6 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B1 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B2 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B4 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C2 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C3 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D1 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D3 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D4 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C3 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C4 = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X13Y132_SLICE_X18Y132_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D2 = CLBLM_R_X5Y124_SLICE_X6Y124_DQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D3 = CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D4 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D5 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D5 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B4 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B5 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C2 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C3 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C4 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A4 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C5 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B4 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B6 = 1'b1;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A1 = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A3 = CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A4 = CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A5 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A6 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C2 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D1 = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B1 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B3 = CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B4 = CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B6 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C2 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C3 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C4 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C5 = CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C6 = CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A1 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A2 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A4 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D2 = CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D2 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D4 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D6 = CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A5 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A6 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B1 = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B2 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A1 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A2 = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A3 = CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A5 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A6 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C1 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D3 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B2 = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B3 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B5 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D2 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C1 = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C3 = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C4 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C5 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A3 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D6 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D4 = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A4 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D6 = CLBLL_L_X4Y123_SLICE_X5Y123_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A6 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A3 = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B2 = CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B3 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B5 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C4 = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C5 = CLBLL_L_X4Y123_SLICE_X4Y123_CQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D1 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D2 = CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D5 = CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A1 = CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A2 = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A3 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A4 = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A5 = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A6 = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B1 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B2 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B6 = CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C1 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C4 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D1 = CLBLL_L_X4Y124_SLICE_X5Y124_C5Q;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D2 = CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D3 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D5 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A1 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A2 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A3 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A5 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A6 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B1 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B2 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B3 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B5 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B6 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C1 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C2 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C3 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C5 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C6 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D1 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D2 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D3 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C5 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D5 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C6 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A1 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A2 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A3 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B1 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B2 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B3 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B5 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C1 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C2 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C3 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C5 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D1 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D2 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D3 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D5 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D6 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A2 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A3 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A5 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A6 = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B1 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B2 = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B3 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B4 = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B5 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B6 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C1 = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C3 = CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C4 = CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C5 = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B1 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B3 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D2 = CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D3 = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D4 = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D6 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_AX = CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A1 = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A2 = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A3 = CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A4 = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A5 = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A6 = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B2 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B3 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B5 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C1 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C2 = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C3 = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C4 = CLBLL_L_X2Y124_SLICE_X0Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C5 = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C6 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D1 = CLBLL_L_X4Y123_SLICE_X4Y123_C5Q;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D4 = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D6 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A2 = CLBLM_L_X10Y128_SLICE_X12Y128_A5Q;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A1 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C6 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D6 = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B2 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B4 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B5 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C1 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C2 = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C3 = CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C4 = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C5 = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C6 = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C5 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D1 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D3 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D5 = CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D6 = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A3 = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A4 = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A6 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C5 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D2 = CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D4 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D5 = CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D6 = CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A1 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A2 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A3 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A4 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D5 = CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B1 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B2 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B3 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B4 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C1 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C2 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C3 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C4 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D1 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D2 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D3 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D4 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A1 = CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A2 = CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A5 = CLBLM_L_X10Y129_SLICE_X13Y129_DQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B1 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B2 = CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B3 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B4 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C1 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C2 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C3 = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C4 = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C5 = CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C6 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D1 = CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D2 = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D3 = CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D4 = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D5 = CLBLM_L_X12Y120_SLICE_X16Y120_BO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D6 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C4 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C5 = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C6 = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B6 = CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D2 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D3 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C4 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D5 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D6 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C6 = CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A5 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B1 = CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B2 = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B3 = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B4 = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B5 = CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B6 = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C1 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C2 = CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C4 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C5 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C6 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D2 = CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D3 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D1 = CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D4 = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D5 = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D6 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B5 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A2 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A3 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A4 = CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A5 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B6 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A6 = CLBLM_R_X3Y128_SLICE_X2Y128_AO5;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B2 = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B4 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B5 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B6 = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C1 = CLBLL_L_X2Y126_SLICE_X1Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C2 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C3 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C4 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C5 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C6 = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B5 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B6 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D1 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D2 = CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D3 = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D4 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D6 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C4 = CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C5 = CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C3 = CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C4 = CLBLM_R_X7Y131_SLICE_X8Y131_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A1 = CLBLM_L_X12Y125_SLICE_X16Y125_DQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A2 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A3 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A5 = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A6 = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C6 = CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B1 = CLBLM_L_X10Y129_SLICE_X13Y129_DQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B2 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B4 = CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B6 = CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C2 = CLBLM_L_X12Y122_SLICE_X17Y122_CQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C4 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C5 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D2 = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D3 = CLBLM_L_X12Y125_SLICE_X16Y125_DQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D4 = CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D6 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A2 = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A3 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A4 = CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A5 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A6 = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B1 = CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B2 = CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B4 = CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B5 = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B6 = CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C1 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C2 = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C3 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C4 = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C5 = CLBLM_R_X3Y128_SLICE_X3Y128_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C6 = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D1 = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D2 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D4 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D5 = CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D6 = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D4 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A1 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A2 = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A3 = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A4 = CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A5 = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A6 = CLBLL_L_X2Y126_SLICE_X0Y126_CO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B1 = CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B2 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B3 = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B4 = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B5 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B6 = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C1 = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C2 = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C3 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C4 = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C5 = CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C6 = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D2 = CLBLM_R_X3Y128_SLICE_X2Y128_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D3 = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D4 = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D5 = CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A1 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A3 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B1 = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B2 = CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B3 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B6 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C1 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C2 = CLBLM_L_X12Y122_SLICE_X17Y122_CQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C5 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C6 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D3 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D4 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D5 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A2 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A5 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A6 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B2 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B6 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C2 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C3 = CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C5 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D1 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D2 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D3 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D4 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D5 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D6 = CLBLM_L_X12Y125_SLICE_X17Y125_CQ;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B1 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B2 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B3 = CLBLM_L_X10Y128_SLICE_X12Y128_DO5;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B6 = CLBLM_R_X3Y128_SLICE_X3Y128_AO5;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C1 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C3 = CLBLM_R_X5Y126_SLICE_X7Y126_CQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C4 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C5 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D2 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D5 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D6 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A4 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B2 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B3 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B4 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B5 = CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C2 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C4 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C5 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C6 = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D1 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D4 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D6 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A1 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A3 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A4 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A5 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B1 = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B3 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B4 = CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B5 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B6 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C1 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C2 = CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C3 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C4 = CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C5 = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C6 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D1 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D2 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D3 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D4 = CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D5 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A1 = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A2 = CLBLM_L_X12Y124_SLICE_X16Y124_BO5;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A3 = CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A4 = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A5 = CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A6 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B1 = CLBLM_L_X12Y124_SLICE_X16Y124_BO5;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B2 = CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B4 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B5 = CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C1 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C2 = CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C3 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C4 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C5 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C6 = CLBLM_L_X12Y125_SLICE_X17Y125_BQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D2 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D3 = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D4 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D5 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D6 = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A1 = CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A3 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A4 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A6 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B2 = CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B3 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B5 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B6 = CLBLL_L_X4Y124_SLICE_X5Y124_CQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C6 = CLBLL_L_X4Y129_SLICE_X4Y129_CQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B2 = CLBLM_R_X5Y128_SLICE_X7Y128_C5Q;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B4 = CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B5 = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C1 = CLBLM_R_X3Y129_SLICE_X2Y129_AO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C4 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C5 = CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C6 = CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D4 = CLBLM_R_X3Y128_SLICE_X3Y128_AO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D5 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D6 = CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A2 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A3 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A6 = CLBLM_L_X12Y124_SLICE_X17Y124_DQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B1 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B2 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B5 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B6 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C1 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C2 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C3 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C5 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D1 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D2 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D3 = CLBLM_L_X12Y124_SLICE_X17Y124_DQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A1 = CLBLM_L_X12Y126_SLICE_X16Y126_A5Q;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A2 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A3 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A4 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A6 = 1'b1;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_AX = CLBLM_R_X11Y123_SLICE_X14Y123_DQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B1 = CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B2 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B3 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B4 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B5 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C1 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C2 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C3 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C4 = CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C5 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D1 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D2 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D3 = CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D4 = CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D5 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D6 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_SR = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D2 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A1 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A2 = CLBLL_L_X4Y129_SLICE_X4Y129_CQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A3 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A5 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_AX = CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B1 = CLBLL_L_X4Y124_SLICE_X5Y124_CQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B2 = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B3 = CLBLM_R_X3Y130_SLICE_X3Y130_CQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B5 = CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C1 = CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C2 = CLBLM_R_X3Y130_SLICE_X3Y130_CQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C4 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C6 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C3 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C4 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C5 = CLBLM_L_X10Y129_SLICE_X13Y129_DQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D2 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D3 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D5 = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C6 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A3 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A4 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A5 = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A1 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A3 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D3 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B2 = CLBLM_L_X12Y125_SLICE_X17Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B4 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B5 = CLBLM_R_X13Y126_SLICE_X18Y126_DQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D5 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C1 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C2 = CLBLM_L_X12Y125_SLICE_X17Y125_CQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C3 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C6 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D6 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D2 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D3 = CLBLM_L_X12Y125_SLICE_X17Y125_DQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D6 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A1 = CLBLM_L_X12Y125_SLICE_X17Y125_DQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A2 = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A3 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A4 = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B1 = CLBLM_L_X12Y124_SLICE_X16Y124_BO5;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B2 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B3 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B4 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B6 = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C1 = CLBLM_L_X12Y124_SLICE_X16Y124_CO5;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C2 = CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C6 = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D1 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D2 = CLBLM_L_X10Y128_SLICE_X12Y128_B5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D3 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D4 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C5 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B4 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B5 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B6 = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C4 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D2 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C5 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A1 = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A3 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A4 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A5 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B1 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B2 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B4 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B5 = CLBLM_R_X3Y131_SLICE_X3Y131_CO5;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C1 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C2 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C3 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C4 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C5 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D1 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D2 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D3 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D4 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D5 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D6 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C6 = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B5 = CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A1 = CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C2 = CLBLM_R_X11Y127_SLICE_X15Y127_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A2 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A3 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A4 = CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C3 = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A6 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B1 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C4 = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C5 = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B6 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C2 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C3 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C4 = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C5 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C6 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D1 = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D2 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D3 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D4 = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D5 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A1 = CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A3 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A4 = CLBLM_L_X12Y126_SLICE_X16Y126_DO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A5 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A6 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C4 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_AX = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C5 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B2 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B3 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B4 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B6 = CLBLM_L_X12Y127_SLICE_X17Y127_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C6 = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C1 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C2 = CLBLM_L_X12Y126_SLICE_X16Y126_CQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C3 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C5 = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C6 = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D1 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D3 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D4 = CLBLM_L_X12Y126_SLICE_X16Y126_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D5 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D2 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D1 = CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A2 = CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A3 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A4 = CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A6 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B2 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B4 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B5 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B6 = CLBLM_R_X13Y126_SLICE_X18Y126_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C1 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C2 = CLBLM_L_X12Y127_SLICE_X17Y127_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C3 = CLBLM_R_X13Y126_SLICE_X18Y126_DQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C5 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C6 = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D1 = CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D2 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D3 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D4 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D5 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A1 = CLBLM_L_X12Y124_SLICE_X17Y124_DQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A2 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A3 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A4 = CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A6 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B1 = CLBLM_R_X11Y127_SLICE_X15Y127_CQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B2 = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B3 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B4 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B6 = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C1 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C3 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C4 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C5 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C6 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D1 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D2 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D3 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D4 = CLBLM_L_X12Y126_SLICE_X16Y126_A5Q;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D5 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D6 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C4 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_R_X11Y123_SLICE_X14Y123_D5Q;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A1 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A2 = CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A3 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A4 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A5 = CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B1 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B2 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B3 = CLBLM_L_X12Y129_SLICE_X17Y129_DO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B4 = CLBLM_R_X13Y126_SLICE_X18Y126_CQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B5 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B6 = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C1 = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C2 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C3 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C4 = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C5 = CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C6 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D1 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D2 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D6 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D4 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D5 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A3 = CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A4 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A5 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A6 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B2 = CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B3 = CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A3 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A6 = CLBLM_L_X8Y121_SLICE_X11Y121_A5Q;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C1 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C2 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B4 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B6 = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D1 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D2 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D3 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C1 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C2 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C4 = CLBLM_L_X8Y121_SLICE_X11Y121_A5Q;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D5 = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D6 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X13Y132_SLICE_X18Y132_AQ;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C2 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A1 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A3 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A4 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A5 = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A6 = CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B1 = CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B2 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B3 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B4 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A1 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C2 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C3 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C4 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C5 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A3 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A4 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A5 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B1 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B5 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D2 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D3 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D4 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C1 = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B3 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B4 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C2 = CLBLM_L_X8Y121_SLICE_X11Y121_A5Q;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D1 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D5 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A2 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A3 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A4 = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A5 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A6 = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D1 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D2 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D4 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D6 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B1 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B3 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B4 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B5 = CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A1 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A2 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A4 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A5 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C1 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C2 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C3 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B3 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B4 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B6 = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D1 = CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D2 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D4 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C1 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D6 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C2 = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D3 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C3 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C4 = CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C6 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C5 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C6 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D2 = CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D3 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D4 = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D5 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D6 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A1 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A2 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A5 = CLBLM_R_X13Y126_SLICE_X18Y126_CQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A6 = CLBLM_L_X12Y122_SLICE_X17Y122_CQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D1 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D2 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B1 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B2 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B4 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B6 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C2 = CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C3 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C4 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C5 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D5 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D6 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D2 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D3 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D5 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D6 = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A2 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A3 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A5 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_DQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B1 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B2 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B3 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C2 = CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C3 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C4 = CLBLM_L_X10Y129_SLICE_X13Y129_DQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C6 = CLBLM_L_X12Y125_SLICE_X17Y125_CQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D1 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D2 = CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D3 = CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D4 = CLBLM_L_X12Y122_SLICE_X17Y122_CQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D5 = CLBLM_L_X12Y125_SLICE_X17Y125_CQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D6 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A6 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C4 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C5 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C6 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B3 = CLBLM_R_X13Y128_SLICE_X19Y128_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B5 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B6 = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C3 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A1 = CLBLM_R_X11Y122_SLICE_X15Y122_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A2 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A3 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A4 = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A5 = CLBLM_L_X10Y128_SLICE_X13Y128_DQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A6 = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B1 = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B2 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B3 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B4 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C1 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C2 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C3 = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C4 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C6 = CLBLM_L_X10Y128_SLICE_X13Y128_D5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D2 = CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D4 = CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D5 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D6 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A1 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A2 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A3 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A4 = CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A5 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_AX = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B2 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B3 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C2 = CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C3 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C4 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_SR = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C5 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C6 = CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B2 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D1 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D3 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D4 = CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D6 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B4 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B4 = CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A3 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B6 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B3 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C3 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D3 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D5 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A2 = CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A3 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A4 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C4 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A6 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C5 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C6 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B3 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C3 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D3 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D5 = CLBLM_L_X10Y128_SLICE_X13Y128_D5Q;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A1 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A3 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C3 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A1 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A3 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A4 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A5 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B1 = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B2 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B6 = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C1 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C2 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C3 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C4 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A3 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_CO5;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D2 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D3 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D4 = CLBLM_L_X10Y121_SLICE_X13Y121_AO5;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D5 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B5 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B6 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D6 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B2 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C1 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C2 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C3 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C4 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C5 = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A1 = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B2 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A6 = CLBLM_L_X10Y127_SLICE_X13Y127_C5Q;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B3 = CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D3 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D4 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D5 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C1 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C2 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C3 = CLBLM_R_X11Y122_SLICE_X15Y122_A5Q;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D2 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D3 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D4 = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D6 = CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A2 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A3 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B2 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B3 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B6 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C2 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C3 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D3 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D4 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D2 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D3 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D6 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D6 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A1 = CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A2 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A4 = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A5 = CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A6 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B2 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B3 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B6 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C2 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D3 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A2 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A6 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_AX = CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B1 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B2 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B6 = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C2 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C3 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C4 = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D1 = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D2 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D4 = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D5 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A1 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A2 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A3 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A6 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B1 = CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B4 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B5 = CLBLM_L_X10Y126_SLICE_X12Y126_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B6 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C3 = CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C5 = CLBLM_L_X10Y126_SLICE_X12Y126_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C6 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D4 = CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D5 = CLBLM_R_X7Y123_SLICE_X8Y123_DQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D6 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A2 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A3 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A5 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B1 = CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B2 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B3 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B4 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B5 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B6 = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C1 = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C4 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C6 = CLBLM_L_X12Y127_SLICE_X17Y127_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D4 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A2 = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A3 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A6 = CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B1 = CLBLM_L_X12Y126_SLICE_X16Y126_CQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B3 = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B4 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B5 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B6 = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C1 = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C2 = CLBLM_R_X13Y126_SLICE_X18Y126_CQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C3 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C4 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C6 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D1 = CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D2 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D3 = CLBLM_R_X13Y126_SLICE_X18Y126_DQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D4 = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D6 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D6 = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A1 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A3 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A4 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A5 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C3 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B1 = CLBLM_R_X11Y123_SLICE_X14Y123_A5Q;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B2 = CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B4 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C2 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C3 = CLBLM_R_X11Y124_SLICE_X15Y124_DQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C4 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D1 = CLBLM_R_X11Y123_SLICE_X14Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D4 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D6 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A2 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A3 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A6 = CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B2 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B3 = CLBLM_R_X11Y123_SLICE_X14Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B4 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B5 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B6 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C1 = CLBLM_L_X10Y123_SLICE_X13Y123_D5Q;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C2 = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C3 = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C4 = CLBLM_L_X10Y128_SLICE_X13Y128_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C5 = CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C6 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D1 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D3 = CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D6 = CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A1 = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A2 = CLBLM_R_X13Y128_SLICE_X19Y128_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A3 = CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A5 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B1 = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B2 = CLBLM_R_X13Y128_SLICE_X19Y128_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B3 = CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B4 = CLBLM_L_X12Y127_SLICE_X17Y127_CQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B5 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B6 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C1 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C2 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C3 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C4 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C5 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C6 = CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D1 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D2 = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D4 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D5 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D6 = CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A1 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A2 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A3 = CLBLM_R_X13Y127_SLICE_X19Y127_AO5;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A4 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A5 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_AX = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B1 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B2 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B3 = CLBLM_R_X13Y127_SLICE_X19Y127_AO5;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B4 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B5 = CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C1 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C2 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C3 = CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C4 = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C5 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C6 = CLBLM_R_X13Y126_SLICE_X18Y126_DQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D1 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D2 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D3 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D4 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D6 = CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_SR = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A1 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A3 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A4 = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_AX = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B1 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B2 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B5 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C3 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C6 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C2 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D6 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D2 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D3 = CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A1 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A4 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B2 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B4 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C4 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C5 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C6 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D3 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D5 = CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D6 = CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D3 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A2 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A3 = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A4 = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A5 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B1 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B2 = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B3 = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B4 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B5 = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B6 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C1 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C2 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C3 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C4 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C5 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C6 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D1 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D2 = CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D3 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D4 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D5 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D6 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A1 = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A2 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A3 = CLBLM_L_X12Y126_SLICE_X16Y126_CQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A4 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D5 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A5 = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A6 = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B1 = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B2 = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B3 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B4 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B5 = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B6 = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C1 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C2 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C3 = CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C4 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C5 = CLBLM_L_X12Y129_SLICE_X17Y129_DO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C6 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D1 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D2 = CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D3 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D4 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D5 = CLBLM_L_X12Y129_SLICE_X17Y129_DO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D6 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C3 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C4 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X3Y130_SLICE_X3Y130_A5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B6 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A1 = CLBLM_L_X10Y125_SLICE_X13Y125_B5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A3 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A4 = CLBLM_L_X12Y125_SLICE_X17Y125_DQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B5 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A1 = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A2 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A4 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C4 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C5 = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C6 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B1 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B2 = CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B4 = CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B6 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C2 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C3 = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C5 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C6 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D6 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D2 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D3 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D4 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A6 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D3 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D4 = CLBLL_L_X4Y121_SLICE_X4Y121_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D5 = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B2 = CLBLM_L_X12Y126_SLICE_X16Y126_A5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B5 = CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C1 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C2 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C3 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C4 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A2 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A3 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A5 = CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D5 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D1 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D2 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B1 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B2 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B3 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B4 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B6 = CLBLL_L_X4Y122_SLICE_X5Y122_AO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C2 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C3 = CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C4 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C5 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D2 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D3 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D4 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D5 = CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A1 = CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A2 = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A4 = CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B4 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A6 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B1 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B5 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B2 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B3 = CLBLM_L_X12Y129_SLICE_X17Y129_DO5;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B4 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B5 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B6 = CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A1 = CLBLM_L_X12Y120_SLICE_X16Y120_AO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A4 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A5 = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A6 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C1 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C2 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C3 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B1 = CLBLM_L_X10Y129_SLICE_X13Y129_DQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B6 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C2 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C3 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C4 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C5 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D3 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D4 = CLBLM_R_X11Y129_SLICE_X15Y129_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A2 = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A3 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A4 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A5 = CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C4 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C4 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B1 = CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A1 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A2 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A4 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A5 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C1 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C2 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C5 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D1 = CLBLM_R_X13Y129_SLICE_X18Y129_CO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D2 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D3 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D4 = CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D5 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D6 = CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D4 = CLBLM_L_X10Y127_SLICE_X13Y127_C5Q;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B2 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B6 = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C1 = CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C2 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A3 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A1 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A2 = CLBLM_R_X7Y122_SLICE_X9Y122_C5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A3 = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A4 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B2 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B3 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A6 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B6 = CLBLM_R_X5Y123_SLICE_X6Y123_DQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B1 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B2 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C1 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C2 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C3 = CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C4 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B3 = CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B4 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B6 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C1 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C2 = CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C3 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C5 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C6 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D6 = CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D2 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D3 = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D1 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D2 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D3 = CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D6 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A3 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A4 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B1 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B2 = CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B4 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B5 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B6 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_BX = CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C1 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C2 = CLBLM_L_X10Y127_SLICE_X13Y127_C5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C3 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C4 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C5 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C6 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A1 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A2 = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A3 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A4 = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B1 = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B2 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B4 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B5 = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D2 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C1 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C2 = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C3 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C4 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C5 = CLBLL_L_X4Y122_SLICE_X5Y122_B5Q;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C6 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D2 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D3 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D4 = CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D5 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D6 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A1 = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A2 = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A3 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A4 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A5 = CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A6 = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B1 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B2 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B3 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B4 = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B5 = CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B6 = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D3 = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C1 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D4 = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C3 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C5 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D5 = CLBLM_R_X11Y127_SLICE_X15Y127_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D6 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D3 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D5 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A1 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A2 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A3 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A4 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A5 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B1 = CLBLM_R_X11Y125_SLICE_X14Y125_DQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B4 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B6 = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C1 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C2 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C3 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C4 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C6 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D2 = CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D5 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D6 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A1 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A2 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A4 = CLBLM_R_X11Y128_SLICE_X15Y128_CQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A6 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A3 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A4 = CLBLM_R_X11Y123_SLICE_X14Y123_D5Q;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A5 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A6 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B6 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B2 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B3 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B5 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B6 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C5 = CLBLM_L_X10Y127_SLICE_X13Y127_C5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C1 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C2 = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C3 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C5 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D1 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D2 = CLBLM_R_X7Y123_SLICE_X8Y123_DQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D6 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D5 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D6 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A3 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A4 = CLBLM_L_X10Y129_SLICE_X13Y129_D5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A5 = CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_AX = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B2 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B6 = CLBLM_R_X7Y127_SLICE_X8Y127_DQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A1 = CLBLL_L_X4Y122_SLICE_X5Y122_B5Q;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A2 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C6 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A3 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A5 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A6 = CLBLM_R_X7Y127_SLICE_X8Y127_D5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C2 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B1 = CLBLL_L_X4Y123_SLICE_X5Y123_CQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B3 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B4 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D2 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B6 = CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D5 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D1 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C2 = CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C4 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C5 = CLBLL_L_X4Y123_SLICE_X5Y123_CQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C6 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D6 = CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D1 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D2 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D3 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D5 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D6 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A2 = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A3 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A5 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B1 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B2 = CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B4 = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B5 = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B6 = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C1 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C2 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C3 = CLBLM_R_X11Y122_SLICE_X15Y122_A5Q;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C4 = CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C5 = CLBLM_R_X11Y124_SLICE_X15Y124_DQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C6 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D1 = CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D2 = CLBLM_L_X12Y125_SLICE_X16Y125_DQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D3 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D4 = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D5 = CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D6 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A1 = CLBLM_R_X11Y121_SLICE_X14Y121_B5Q;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A3 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B2 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B3 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B4 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C1 = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C2 = CLBLM_L_X12Y121_SLICE_X16Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C3 = CLBLM_L_X10Y128_SLICE_X13Y128_DQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C5 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C6 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D3 = CLBLM_R_X11Y123_SLICE_X14Y123_A5Q;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D4 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D5 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D6 = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A1 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A2 = CLBLM_R_X7Y122_SLICE_X9Y122_C5Q;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A3 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A4 = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A3 = CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A4 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A5 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B1 = CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B3 = CLBLM_L_X10Y128_SLICE_X13Y128_CQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B6 = CLBLM_L_X10Y129_SLICE_X12Y129_CQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C4 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C5 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D1 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D2 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D1 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D5 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A1 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A2 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_AX = CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B2 = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B3 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A1 = CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A2 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_BX = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C2 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C3 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B2 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B3 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C5 = CLBLM_R_X11Y129_SLICE_X15Y129_CQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D1 = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C2 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C3 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C5 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D2 = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D3 = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D1 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D6 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A3 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A4 = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A5 = CLBLM_R_X11Y128_SLICE_X15Y128_DQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A6 = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_AX = CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D4 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B1 = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B2 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B3 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B4 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B6 = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A4 = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C1 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C4 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C6 = CLBLM_L_X12Y125_SLICE_X17Y125_BQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D4 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A2 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A3 = CLBLM_R_X13Y132_SLICE_X18Y132_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A4 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D4 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D5 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D6 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A1 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A2 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A4 = CLBLM_R_X11Y121_SLICE_X14Y121_B5Q;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B1 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B2 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B3 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B5 = CLBLM_R_X7Y130_SLICE_X8Y130_A5Q;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C1 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A6 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C2 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C4 = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A4 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C5 = CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C6 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A5 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D2 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D3 = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D4 = CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D5 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B3 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_D5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B5 = CLBLL_L_X4Y123_SLICE_X4Y123_C5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C1 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C2 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C3 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A1 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A2 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C4 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A3 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A4 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A6 = CLBLL_L_X4Y127_SLICE_X4Y127_A5Q;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C5 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B1 = CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A5 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B2 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B3 = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B4 = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B5 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B6 = CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B2 = CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B4 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B5 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C1 = CLBLL_L_X4Y127_SLICE_X4Y127_CO5;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C1 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C2 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C4 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C5 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D1 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D2 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D3 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D4 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A1 = CLBLM_L_X10Y130_SLICE_X12Y130_A5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A2 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A5 = CLBLM_R_X11Y129_SLICE_X15Y129_CQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D2 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B2 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B3 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B5 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D3 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C4 = CLBLM_L_X10Y127_SLICE_X12Y127_AO5;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C6 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C2 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C1 = CLBLL_L_X4Y127_SLICE_X4Y127_CO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C2 = CLBLL_L_X4Y122_SLICE_X5Y122_B5Q;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C3 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C4 = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C5 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C3 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D1 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D2 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D3 = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D4 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D5 = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D6 = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A1 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A3 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A4 = CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A5 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B2 = CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B3 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B4 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B5 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C3 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C2 = CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C3 = CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C6 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D1 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D2 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D3 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D4 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D5 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A1 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A3 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A4 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A5 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A6 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B2 = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B4 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B5 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C1 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C3 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C5 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D3 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D5 = CLBLM_L_X8Y124_SLICE_X10Y124_C5Q;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D6 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X10Y123_SLICE_X13Y123_DQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A4 = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D5 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A5 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B4 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B5 = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A1 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A2 = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A3 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A4 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A5 = CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A6 = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B1 = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B2 = CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B3 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B4 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B5 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B6 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A2 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A6 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C1 = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C3 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C4 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C6 = CLBLM_R_X5Y122_SLICE_X7Y122_DQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B1 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B2 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B3 = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B4 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B5 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B6 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A1 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D1 = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D3 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D5 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D6 = CLBLL_L_X4Y127_SLICE_X4Y127_DO5;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A3 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B6 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B1 = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B2 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C2 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C4 = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C5 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D3 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D4 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A2 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A3 = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A1 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A3 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A4 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A5 = CLBLM_L_X8Y128_SLICE_X10Y128_B5Q;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D2 = CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D3 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A4 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A2 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B2 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C1 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C2 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C5 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D3 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D4 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D5 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D2 = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A6 = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B1 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C1 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C2 = CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A1 = CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B1 = CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B4 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B5 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C3 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D4 = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D6 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A3 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A4 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A5 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A6 = CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B2 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B4 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C1 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C2 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C4 = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X11Y123_SLICE_X14Y123_DQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D2 = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D3 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D1 = CLBLM_R_X11Y123_SLICE_X15Y123_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D2 = CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D3 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D4 = CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D5 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D6 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B6 = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A2 = CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A3 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A4 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B1 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B2 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B3 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B5 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B6 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A6 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A1 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A3 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A5 = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B1 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B2 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A1 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A2 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A3 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A5 = CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B1 = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B2 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B3 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B5 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B6 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D2 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C1 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C2 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C4 = CLBLM_L_X8Y121_SLICE_X11Y121_A5Q;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C5 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C6 = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D4 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A2 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A1 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A3 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A4 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A5 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A6 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D6 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B1 = CLBLL_L_X4Y128_SLICE_X5Y128_B5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B2 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B3 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B5 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A2 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A3 = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A5 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B2 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B3 = CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B5 = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C2 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C3 = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C4 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C5 = CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D5 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D2 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D3 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D4 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D6 = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A1 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_D5Q;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A4 = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B1 = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B2 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B4 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B5 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C2 = CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C4 = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C5 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D4 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D1 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D4 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D5 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A6 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A2 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A3 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A4 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B1 = CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B2 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B4 = CLBLM_R_X11Y123_SLICE_X15Y123_CQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B6 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C4 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C5 = CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C6 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D2 = CLBLM_L_X8Y124_SLICE_X10Y124_C5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D3 = CLBLM_R_X11Y125_SLICE_X14Y125_DQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D4 = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C4 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C5 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A2 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A3 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A4 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A5 = CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A6 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_AX = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B1 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B2 = CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B3 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B5 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C1 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C5 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A1 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A3 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A4 = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A5 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A6 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D1 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D2 = CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D3 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D4 = CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D5 = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A2 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A3 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A6 = CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_AX = CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B3 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B4 = CLBLM_L_X10Y129_SLICE_X12Y129_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C2 = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C3 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C4 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A1 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A2 = CLBLM_R_X3Y130_SLICE_X3Y130_CQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A3 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A6 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B2 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B4 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B5 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D4 = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D6 = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A1 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C4 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C5 = CLBLL_L_X4Y127_SLICE_X4Y127_A5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C6 = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A6 = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D3 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D4 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D5 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D6 = CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C2 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C3 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C6 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D2 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D3 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D5 = CLBLM_R_X11Y123_SLICE_X14Y123_A5Q;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D6 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A3 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A4 = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A5 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B1 = CLBLM_R_X11Y124_SLICE_X15Y124_DQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B2 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B4 = CLBLM_L_X12Y126_SLICE_X16Y126_CQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C2 = CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C4 = CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C5 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C6 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B2 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D3 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D6 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_DQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B5 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A3 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A4 = CLBLM_L_X12Y127_SLICE_X17Y127_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B2 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B3 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B4 = CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B5 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C1 = CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C3 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C4 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C5 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D1 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D2 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D3 = CLBLM_R_X11Y126_SLICE_X14Y126_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D4 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D5 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D6 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A1 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A2 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A3 = CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A4 = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A6 = CLBLM_R_X3Y130_SLICE_X3Y130_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B1 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B2 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B5 = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C1 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C2 = CLBLL_L_X4Y129_SLICE_X4Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C4 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C5 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D1 = CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D4 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A4 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A6 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B1 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B2 = CLBLM_L_X12Y125_SLICE_X16Y125_DQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B3 = CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B4 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B5 = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B6 = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C1 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A3 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A4 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A5 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C2 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C3 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B1 = CLBLL_L_X4Y124_SLICE_X5Y124_CQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B2 = CLBLL_L_X4Y128_SLICE_X5Y128_B5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B3 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B4 = CLBLM_L_X8Y128_SLICE_X10Y128_B5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B6 = CLBLL_L_X4Y129_SLICE_X4Y129_B5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_D5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D2 = CLBLM_L_X10Y123_SLICE_X13Y123_C5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C2 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C3 = CLBLM_L_X8Y128_SLICE_X10Y128_B5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C5 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D6 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A1 = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A3 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A4 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A5 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C6 = CLBLL_L_X4Y127_SLICE_X4Y127_A5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D2 = CLBLL_L_X4Y128_SLICE_X5Y128_B5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D4 = CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D5 = CLBLL_L_X4Y124_SLICE_X5Y124_CQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D6 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B2 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B4 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C4 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C3 = CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C6 = 1'b1;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D3 = CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D4 = CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D5 = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A1 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A3 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A4 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A5 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A6 = CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B2 = CLBLM_R_X11Y127_SLICE_X15Y127_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B4 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B5 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C1 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C2 = CLBLM_R_X11Y127_SLICE_X15Y127_CQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C3 = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D2 = CLBLM_R_X11Y127_SLICE_X15Y127_CQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D3 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D4 = CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D5 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A1 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A2 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A3 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A5 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A6 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B1 = CLBLM_L_X12Y121_SLICE_X16Y121_CQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B2 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B3 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C1 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C2 = CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C3 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C6 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D2 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D3 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D4 = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D6 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A2 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A3 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A5 = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A6 = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C2 = CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B1 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B2 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B4 = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B5 = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B6 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C4 = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C1 = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C2 = CLBLL_L_X4Y130_SLICE_X4Y130_CQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C4 = CLBLM_R_X7Y130_SLICE_X8Y130_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C5 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C6 = CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C6 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D1 = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D2 = CLBLM_R_X3Y130_SLICE_X3Y130_DO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D3 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D5 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D6 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A1 = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A2 = CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A3 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A4 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A5 = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B2 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B3 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B5 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A2 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A3 = CLBLM_R_X7Y130_SLICE_X8Y130_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A4 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C1 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C3 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C4 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C5 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A5 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A6 = CLBLL_L_X4Y130_SLICE_X4Y130_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_AX = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B1 = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B3 = CLBLM_L_X8Y128_SLICE_X10Y128_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B4 = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B5 = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B6 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C1 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C2 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C4 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C3 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C6 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C5 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A3 = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A4 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D1 = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D3 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D4 = CLBLL_L_X4Y124_SLICE_X5Y124_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B3 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D5 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D6 = CLBLL_L_X4Y127_SLICE_X4Y127_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B6 = CLBLM_L_X8Y124_SLICE_X10Y124_AO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B4 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B5 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C1 = CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C2 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C4 = CLBLM_L_X10Y123_SLICE_X13Y123_C5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C4 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D6 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C5 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D1 = CLBLM_R_X7Y123_SLICE_X9Y123_AO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D2 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D3 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D4 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D5 = CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D6 = CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C6 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C2 = CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A2 = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A6 = CLBLM_L_X10Y128_SLICE_X12Y128_B5Q;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C4 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_AX = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C5 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B2 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B4 = CLBLM_R_X11Y128_SLICE_X15Y128_DQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B5 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C1 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C2 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C5 = CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D3 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D5 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D2 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D4 = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D5 = CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D6 = CLBLM_R_X11Y128_SLICE_X15Y128_DQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A1 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A2 = CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A3 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_AX = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B3 = CLBLM_L_X12Y125_SLICE_X17Y125_CQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B4 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B5 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B6 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A1 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C2 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A2 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C4 = CLBLM_R_X11Y128_SLICE_X14Y128_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C6 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A4 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D2 = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A5 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D3 = CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D4 = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D5 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D6 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A3 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A4 = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A5 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A6 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_AX = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B5 = CLBLM_L_X12Y125_SLICE_X16Y125_D5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B3 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B4 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B5 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C2 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C3 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C4 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C5 = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D6 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A2 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A3 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A4 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C6 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B1 = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C2 = CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C1 = CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C3 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D1 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D4 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D5 = CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D6 = CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A1 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A4 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A5 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B1 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B3 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B4 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B5 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C2 = CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C3 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C4 = CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C5 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C6 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D1 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D2 = CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D3 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D4 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D5 = CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D6 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D5 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A1 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A2 = CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A3 = CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B1 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B3 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B4 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B5 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A5 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A6 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C1 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C2 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C3 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D3 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D4 = CLBLM_R_X11Y125_SLICE_X14Y125_DQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A1 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A2 = CLBLM_L_X10Y129_SLICE_X12Y129_CQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A3 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A5 = CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B3 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A2 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A4 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A6 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C2 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C3 = CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B2 = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B3 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B4 = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B5 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D1 = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D4 = CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C1 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C3 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C4 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C5 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C6 = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D5 = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D2 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D5 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A1 = CLBLM_R_X11Y129_SLICE_X14Y129_CQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A2 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A3 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A6 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B1 = CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B5 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B6 = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A1 = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A2 = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A4 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C1 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C6 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D2 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D4 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D6 = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A1 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A3 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_AX = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B1 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B3 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B4 = CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B5 = CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B6 = CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C1 = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C3 = CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C4 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C6 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D4 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D6 = CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D1 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D2 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_SR = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A3 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A5 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A6 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A3 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A4 = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C2 = CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_AX = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B2 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B4 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B6 = CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C2 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C3 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5 = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C6 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A2 = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A4 = CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D2 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D3 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D4 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B3 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A2 = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A3 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A4 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A5 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C2 = CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_AX = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B2 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B5 = CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D2 = CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C2 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C3 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C6 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D5 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D2 = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D3 = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D4 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A4 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B2 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B4 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B5 = CLBLM_R_X11Y128_SLICE_X15Y128_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C2 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C3 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C4 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C5 = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D2 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D3 = CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A2 = CLBLM_L_X10Y128_SLICE_X13Y128_D5Q;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A4 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A6 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B1 = CLBLM_L_X10Y128_SLICE_X12Y128_A5Q;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B2 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B4 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B6 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C2 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C5 = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C6 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D2 = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D4 = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X13Y132_SLICE_X18Y132_AQ;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A1 = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A2 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A3 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A4 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A5 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A6 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B1 = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B2 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B3 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B4 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B5 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B6 = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = CLBLM_R_X5Y126_SLICE_X7Y126_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C1 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C2 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C3 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D1 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A1 = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A2 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A3 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A4 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A6 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B2 = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B3 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C1 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C2 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C3 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D2 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = CLBLL_L_X4Y129_SLICE_X4Y129_B5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D3 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D4 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D6 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_DQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D5 = CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A1 = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A6 = CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B4 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C5 = CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C6 = CLBLM_L_X10Y123_SLICE_X13Y123_D5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D2 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D3 = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D4 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D5 = CLBLM_L_X10Y128_SLICE_X12Y128_A5Q;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A2 = CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A6 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B1 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B2 = CLBLM_R_X7Y130_SLICE_X8Y130_A5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B3 = CLBLM_R_X11Y129_SLICE_X14Y129_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A6 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C2 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C4 = CLBLM_R_X11Y129_SLICE_X14Y129_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C5 = CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C6 = CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D1 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D4 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B4 = CLBLM_R_X5Y121_SLICE_X7Y121_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A2 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A3 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A4 = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A6 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C4 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B1 = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B2 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B4 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C1 = CLBLM_R_X7Y122_SLICE_X9Y122_C5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C2 = CLBLM_L_X10Y123_SLICE_X13Y123_D5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C4 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D3 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D4 = CLBLM_L_X10Y128_SLICE_X13Y128_D5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D5 = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D6 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_AX = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A1 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A2 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A4 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B2 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B3 = CLBLM_R_X5Y122_SLICE_X6Y122_DQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B6 = CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C1 = CLBLM_L_X12Y125_SLICE_X16Y125_D5Q;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C2 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C4 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C6 = CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_SR = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D2 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D6 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X3Y130_SLICE_X3Y130_CQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_R_X11Y123_SLICE_X14Y123_D5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A1 = CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A2 = CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A3 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A4 = CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A5 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A6 = CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B1 = CLBLM_L_X10Y129_SLICE_X12Y129_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B2 = CLBLM_R_X11Y129_SLICE_X14Y129_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B3 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B4 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B5 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B6 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C1 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C4 = CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C6 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D1 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D2 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D6 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A2 = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A5 = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B2 = CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B4 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B5 = CLBLM_L_X8Y123_SLICE_X10Y123_CO5;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C1 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C2 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C3 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D1 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D2 = CLBLM_R_X11Y128_SLICE_X15Y128_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D4 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D5 = CLBLM_L_X10Y123_SLICE_X13Y123_D5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D6 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C2 = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C3 = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C5 = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A1 = CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A3 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A4 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D6 = CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A5 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B1 = CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B2 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B3 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B5 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C1 = CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C2 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C3 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C4 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C5 = CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D1 = CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D1 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D2 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D2 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D3 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D4 = CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D5 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D6 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A1 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A2 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A4 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A6 = 1'b1;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B1 = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B2 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B4 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B6 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C3 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C4 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C5 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B1 = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D2 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D4 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D5 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D6 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D3 = CLBLM_R_X7Y123_SLICE_X8Y123_DQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B3 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B5 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B6 = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C1 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A3 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A4 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A1 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A2 = CLBLM_L_X10Y123_SLICE_X13Y123_DQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A3 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A4 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A6 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A5 = CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B1 = CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B4 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B5 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C2 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C3 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C5 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D1 = CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D2 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D3 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D4 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D5 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D1 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D2 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A2 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D3 = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D4 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A4 = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A2 = CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B1 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B2 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B3 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B4 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B6 = CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D5 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D6 = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A2 = CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C2 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C3 = CLBLM_L_X8Y128_SLICE_X10Y128_B5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C4 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C5 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C6 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A3 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A5 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B5 = CLBLL_L_X2Y123_SLICE_X1Y123_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B6 = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_AX = CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B2 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B3 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D2 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D4 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D5 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C1 = CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C2 = CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C4 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C5 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D1 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D2 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D5 = CLBLM_R_X5Y122_SLICE_X6Y122_DQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D6 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A2 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B2 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B4 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A1 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A4 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A5 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C2 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B2 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B4 = CLBLM_R_X7Y123_SLICE_X9Y123_AO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B5 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C1 = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C2 = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C4 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D4 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A3 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A4 = CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D2 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D3 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D4 = CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D5 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B2 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B4 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A4 = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A5 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B1 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B2 = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B4 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C4 = CLBLM_L_X10Y128_SLICE_X13Y128_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C6 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D4 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D1 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D2 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D3 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D5 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D6 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X11Y123_SLICE_X14Y123_DQ;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A2 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A3 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A5 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A6 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_AX = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B1 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B3 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B4 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B5 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C1 = CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C2 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C6 = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C5 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C6 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D1 = CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D3 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D4 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D5 = CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D6 = CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A1 = CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A4 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A5 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A6 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B1 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B2 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A1 = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A3 = CLBLL_L_X2Y123_SLICE_X1Y123_AQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A6 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B4 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B5 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B4 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B5 = CLBLL_L_X4Y123_SLICE_X4Y123_C5Q;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C1 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C1 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C2 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C3 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C4 = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D1 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D5 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C5 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C6 = CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D2 = CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D3 = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D4 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D5 = CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D6 = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A1 = CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A2 = CLBLM_L_X10Y128_SLICE_X13Y128_DQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A3 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A6 = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B2 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B4 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B6 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C1 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C2 = CLBLM_R_X5Y124_SLICE_X6Y124_DQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D2 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C3 = CLBLM_R_X5Y123_SLICE_X6Y123_DQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C4 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C5 = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C6 = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D3 = CLBLM_L_X10Y129_SLICE_X12Y129_DQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D4 = CLBLM_R_X7Y127_SLICE_X8Y127_DQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D1 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D2 = CLBLM_L_X10Y128_SLICE_X13Y128_DQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D3 = CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A2 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A3 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A4 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A6 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B2 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B4 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B5 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B6 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C2 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C3 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C6 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B6 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D1 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D2 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D4 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D5 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D6 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C3 = 1'b1;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C4 = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X3Y130_SLICE_X3Y130_A5Q;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A5 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A6 = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B2 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A5 = CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A6 = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B6 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C4 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_AX = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C3 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D4 = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D6 = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D3 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D5 = CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_SR = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A1 = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A2 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A3 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A4 = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A1 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A3 = CLBLL_L_X2Y123_SLICE_X1Y123_AQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A4 = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A5 = CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A6 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B1 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B3 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B1 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B2 = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B4 = CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B6 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C1 = CLBLL_L_X2Y123_SLICE_X1Y123_AQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C2 = CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C4 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C5 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C6 = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C5 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D4 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D1 = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D2 = CLBLL_L_X2Y126_SLICE_X1Y126_CO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D3 = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D4 = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D5 = CLBLL_L_X2Y125_SLICE_X0Y125_BO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D6 = CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A1 = CLBLL_L_X4Y128_SLICE_X5Y128_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A2 = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A3 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A5 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_AX = CLBLM_R_X7Y126_SLICE_X9Y126_CO5;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B1 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B4 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B5 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C1 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C2 = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C4 = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D3 = CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D4 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D5 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X10Y123_SLICE_X13Y123_DQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A1 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A2 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A4 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A6 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B1 = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B5 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B6 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C1 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C2 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C3 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C4 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D1 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D2 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D4 = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B1 = CLBLM_R_X13Y123_SLICE_X19Y123_CQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A3 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D2 = CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C4 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C5 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D4 = CLBLM_R_X11Y122_SLICE_X15Y122_A5Q;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D2 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D4 = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D5 = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A1 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B1 = CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B2 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B3 = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B4 = CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B5 = CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B6 = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C1 = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C2 = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C3 = CLBLL_L_X2Y125_SLICE_X0Y125_BO5;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C4 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C5 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C6 = CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A4 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A5 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D2 = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D4 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D5 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D6 = CLBLL_L_X2Y124_SLICE_X1Y124_BO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A3 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A4 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A5 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A6 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B1 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B5 = CLBLM_L_X10Y123_SLICE_X13Y123_D5Q;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C2 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C3 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D1 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D2 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D3 = CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D4 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D5 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A2 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A5 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B3 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B4 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B6 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C2 = CLBLM_L_X8Y129_SLICE_X10Y129_DO5;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C4 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D2 = CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D3 = CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A6 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B1 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B2 = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B3 = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B4 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B5 = CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B6 = CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A3 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C1 = CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C2 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C3 = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C4 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A3 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A5 = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A6 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C5 = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C6 = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B4 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D1 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D2 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D3 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D5 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D6 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D6 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A1 = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A6 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A3 = CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A4 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A6 = CLBLM_R_X5Y126_SLICE_X6Y126_DQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B6 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B1 = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B2 = CLBLL_L_X2Y126_SLICE_X0Y126_BO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B3 = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B5 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C6 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C2 = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C3 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C4 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C5 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C6 = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D1 = CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D2 = CLBLL_L_X2Y128_SLICE_X1Y128_CO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D3 = CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D4 = CLBLL_L_X2Y126_SLICE_X1Y126_CO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D5 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D6 = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D2 = 1'b1;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A3 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A4 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A5 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A6 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B2 = CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B4 = CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B5 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C2 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_DQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C6 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D1 = CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D2 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D3 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D4 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D6 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A3 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A4 = CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A6 = CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B1 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B2 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B3 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B6 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C1 = CLBLM_L_X10Y128_SLICE_X12Y128_A5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C2 = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C3 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B2 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C5 = CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C6 = CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D2 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D4 = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D6 = CLBLM_R_X7Y126_SLICE_X9Y126_A5Q;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C4 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A2 = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A4 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A5 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A6 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B5 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B6 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C2 = CLBLM_L_X8Y127_SLICE_X11Y127_B5Q;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C3 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C4 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C6 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A2 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D1 = CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_AX = CLBLM_L_X12Y135_SLICE_X16Y135_AO5;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D2 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D3 = CLBLL_L_X2Y126_SLICE_X0Y126_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D4 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D5 = CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D6 = CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C2 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D2 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A1 = CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A2 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A3 = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A4 = CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A5 = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A6 = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A2 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B2 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B2 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C2 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C3 = CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A3 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D3 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C2 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A5 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D1 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D2 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D3 = CLBLM_R_X3Y128_SLICE_X2Y128_AO5;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D4 = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D5 = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D6 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D2 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A1 = CLBLM_R_X3Y130_SLICE_X3Y130_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A3 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A4 = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_AX = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C1 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B1 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B2 = CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B3 = CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C2 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C3 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C1 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C2 = CLBLM_L_X10Y123_SLICE_X13Y123_D5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C4 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C5 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C5 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C6 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D1 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D2 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D4 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D5 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B4 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A2 = CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B5 = CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A3 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A6 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B6 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_AX = CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B3 = CLBLM_R_X7Y127_SLICE_X8Y127_D5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B4 = CLBLM_R_X7Y131_SLICE_X8Y131_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C2 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C4 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D3 = CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D4 = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D2 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D5 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C4 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D5 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C5 = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D6 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B1 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B2 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B3 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B4 = CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B6 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C6 = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D2 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D5 = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D6 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_AX = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B2 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B1 = CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B3 = CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B2 = CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B3 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B4 = CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B5 = CLBLM_R_X3Y128_SLICE_X2Y128_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B6 = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C1 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C2 = CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C3 = CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C4 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C5 = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C6 = CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B6 = CLBLM_R_X11Y128_SLICE_X14Y128_A5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B5 = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D2 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D3 = CLBLL_L_X2Y129_SLICE_X1Y129_AO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D5 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C3 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C4 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C5 = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C6 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A1 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A2 = CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A3 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A6 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C4 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B1 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B4 = CLBLM_R_X11Y126_SLICE_X14Y126_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B5 = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A1 = CLBLM_R_X7Y120_SLICE_X8Y120_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A4 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C2 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B1 = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B2 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B4 = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B6 = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D3 = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C2 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D4 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C3 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C4 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5 = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C6 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D5 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A2 = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D6 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D2 = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D3 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D4 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B2 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B4 = CLBLM_R_X7Y127_SLICE_X8Y127_DQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B5 = CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B6 = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B1 = CLBLL_L_X4Y130_SLICE_X4Y130_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A2 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A3 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C1 = CLBLM_R_X7Y130_SLICE_X8Y130_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C2 = CLBLM_L_X12Y125_SLICE_X17Y125_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B2 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B4 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B3 = CLBLL_L_X4Y127_SLICE_X4Y127_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B6 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B5 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C1 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C4 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D2 = CLBLM_R_X7Y127_SLICE_X8Y127_DQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D3 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D6 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D1 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D5 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B5 = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B6 = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C5 = CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A1 = CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A3 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A6 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B1 = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B2 = CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B4 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B5 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B6 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A2 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A3 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A6 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C1 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C2 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C3 = CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B2 = CLBLM_R_X5Y121_SLICE_X7Y121_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B5 = CLBLL_L_X4Y121_SLICE_X4Y121_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B6 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D1 = CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C1 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C2 = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C5 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B2 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C6 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D4 = CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A1 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A2 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A3 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A4 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D1 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D4 = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D5 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D6 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A6 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C4 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B1 = CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B2 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A1 = CLBLL_L_X4Y122_SLICE_X5Y122_AO5;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A2 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A3 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A6 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C5 = CLBLM_R_X7Y130_SLICE_X8Y130_A5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B1 = CLBLL_L_X4Y122_SLICE_X5Y122_B5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B2 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D1 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C1 = CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C2 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C3 = CLBLM_L_X12Y121_SLICE_X16Y121_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D5 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D6 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D1 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D2 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B4 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D2 = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D5 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D6 = CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D2 = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D5 = CLBLM_L_X12Y125_SLICE_X16Y125_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A2 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A3 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A4 = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B2 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B4 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B6 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C3 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A3 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A4 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B1 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C6 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B2 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B3 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B4 = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B5 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A1 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A3 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A5 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A6 = CLBLL_L_X4Y123_SLICE_X4Y123_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B1 = CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B2 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B6 = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C1 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C3 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C4 = CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C5 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C6 = CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A4 = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D2 = CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D3 = CLBLM_R_X5Y122_SLICE_X7Y122_DQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D5 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A6 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B1 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B2 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B3 = CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B4 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A1 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A3 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A4 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A6 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C1 = CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C2 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B1 = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B3 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D4 = CLBLL_L_X4Y128_SLICE_X5Y128_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C4 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D2 = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D3 = CLBLM_R_X5Y122_SLICE_X6Y122_DQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D4 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D6 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D6 = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A1 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A2 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A3 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A5 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A6 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B3 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B4 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B5 = CLBLM_R_X7Y126_SLICE_X8Y126_D5Q;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B6 = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C2 = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C5 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C6 = CLBLM_R_X5Y121_SLICE_X7Y121_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D2 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D4 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D5 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D6 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A2 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A3 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A4 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A5 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A6 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B6 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B1 = CLBLM_L_X10Y124_SLICE_X12Y124_DQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B2 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B3 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B5 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B6 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C1 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C2 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C3 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C4 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C1 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D2 = CLBLL_L_X4Y124_SLICE_X5Y124_C5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C2 = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D4 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D5 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C3 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C1 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D2 = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A2 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B4 = CLBLL_L_X2Y128_SLICE_X1Y128_BO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B6 = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C1 = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B3 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B4 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B5 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B6 = CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B4 = CLBLM_R_X5Y123_SLICE_X6Y123_DQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C1 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A1 = CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A2 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A3 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A5 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A6 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C3 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B1 = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B2 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B3 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B4 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B5 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C4 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C5 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C1 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C3 = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C6 = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C5 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C6 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D1 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D2 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D3 = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D4 = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D5 = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B6 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A1 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A4 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A6 = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B2 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B4 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B6 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C4 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C6 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D1 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D3 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D5 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C4 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D5 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C5 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D6 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C6 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A1 = CLBLM_L_X10Y125_SLICE_X13Y125_B5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLM_R_X37Y122_SLICE_X56Y122_AO6;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A4 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A5 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A6 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D5 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B6 = 1'b1;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B1 = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B3 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B5 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B6 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C1 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C2 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D5 = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C5 = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C6 = CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D6 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A1 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A2 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A3 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A4 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A6 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C4 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B1 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B2 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B3 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B4 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B5 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B6 = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C1 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C2 = CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D2 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C4 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C5 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C6 = CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D3 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X3Y130_SLICE_X3Y130_CQ;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D4 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C5 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D1 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D2 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D3 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D4 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D6 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D6 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A1 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A2 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A6 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B1 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B2 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B5 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B6 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C2 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C3 = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C4 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C5 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C6 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D2 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D4 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D6 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A2 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A3 = CLBLM_R_X13Y132_SLICE_X18Y132_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A4 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C5 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C3 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C4 = CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C5 = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X3Y130_SLICE_X3Y130_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A1 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A2 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A4 = CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_AX = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B1 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B2 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B4 = CLBLM_R_X5Y122_SLICE_X7Y122_DQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C6 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C2 = CLBLM_R_X5Y126_SLICE_X7Y126_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C4 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C5 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C6 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D2 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D3 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D4 = CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D5 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A1 = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A2 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A4 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C4 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A3 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B2 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B4 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B5 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B6 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A5 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C5 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C6 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C1 = CLBLM_R_X5Y123_SLICE_X6Y123_DQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C2 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C4 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C5 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D1 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D2 = CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D3 = CLBLM_R_X5Y126_SLICE_X6Y126_DQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C5 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C6 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B5 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B6 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D5 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D6 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B5 = CLBLM_R_X7Y126_SLICE_X9Y126_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C5 = 1'b1;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C5 = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A2 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A4 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A5 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A6 = CLBLM_R_X11Y127_SLICE_X15Y127_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C6 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B2 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B4 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B5 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B6 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C3 = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C5 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C6 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A3 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A4 = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A5 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D1 = CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D2 = CLBLL_L_X4Y127_SLICE_X4Y127_DO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D3 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D4 = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D5 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A1 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A2 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A4 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B1 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B3 = CLBLM_L_X12Y122_SLICE_X16Y122_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B4 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B6 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C2 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C4 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C5 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C6 = CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D2 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D3 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D4 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D4 = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D5 = CLBLM_R_X5Y124_SLICE_X7Y124_CO5;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A2 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A3 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A5 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A6 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B2 = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B5 = CLBLM_R_X5Y128_SLICE_X7Y128_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C1 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C2 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C3 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C5 = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A1 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A2 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A4 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A5 = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_DQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B3 = CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B5 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C1 = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C1 = CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C2 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C3 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C4 = CLBLM_L_X10Y128_SLICE_X12Y128_CO5;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C6 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C4 = CLBLL_L_X4Y129_SLICE_X4Y129_B5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D1 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D2 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B4 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
endmodule
