module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5Q;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CLK;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CLK;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5Q;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5Q;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CLK;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5Q;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CLK;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CLK;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CLK;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5Q;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CLK;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CLK;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BQ;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CLK;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CQ;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CMUX;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AQ;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CLK;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BQ;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CLK;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CQ;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AQ;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BQ;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CLK;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AQ;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CLK;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CLK;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AQ;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BQ;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CLK;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CLK;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CLK;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CLK;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D5Q;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B5Q;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CLK;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D5Q;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CLK;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CLK;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CLK;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CLK;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CLK;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5Q;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C5Q;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CLK;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C5Q;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CLK;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D5Q;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CLK;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C5Q;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D5Q;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C5Q;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CE;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_SR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CLK;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DMUX;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AQ;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CLK;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AQ;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CLK;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BMUX;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CLK;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CMUX;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DMUX;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CLK;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D5Q;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DMUX;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CLK;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B5Q;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BMUX;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CLK;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_DO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_AO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_AO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_BO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_BO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CLK;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CMUX;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_DO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_DO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A5Q;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CLK;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_DMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_DO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_DO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CLK;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_DMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CLK;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_DO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_DQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CLK;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_DO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CLK;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_DQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_AO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_AO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_BO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_BO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CLK;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_DO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_DO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AMUX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CE;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CLK;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DMUX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_SR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DMUX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BMUX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CLK;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CMUX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_DO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CLK;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CMUX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_DO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BMUX;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CLK;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CMUX;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CLK;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_DO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AMUX;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AX;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CE;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CLK;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_DO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_SR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AMUX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CLK;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CQ;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CLK;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CLK;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CLK;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DMUX;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CLK;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CLK;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5Q;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CLK;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CLK;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CLK;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5Q;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CLK;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AQ;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BQ;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CLK;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CLK;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CLK;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5Q;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CLK;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CLK;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CLK;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CMUX;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D5Q;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DMUX;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CLK;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B5Q;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CLK;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AMUX;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AMUX;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AMUX;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AQ;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BQ;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CLK;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AQ;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CLK;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AQ;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CLK;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A5Q;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AQ;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CLK;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CQ;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A5Q;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CLK;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A5Q;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CLK;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AQ;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CLK;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A5Q;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CLK;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CLK;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AMUX;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BMUX;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CLK;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DMUX;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CLK;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CLK;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CE;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CLK;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_SR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CLK;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B5Q;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CLK;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CLK;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C5Q;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A5Q;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CLK;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CLK;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A5Q;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AMUX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AX;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_BO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CLK;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_DO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_BO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_CO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_CO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_DO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_DO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_AO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_AQ;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_BO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_BQ;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CLK;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CQ;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_DO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_DQ;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_AO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_BO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_BO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_CO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_CO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_DO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_DO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_BO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_BO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CLK;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_AO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_BO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_CO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_DO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_DO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_AO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_AO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_BO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_BQ;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_CLK;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_CO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_CQ;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_DMUX;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_DO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_AO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_AQ;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_BO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_BO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_BQ;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_CLK;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_CO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_CO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_DO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_DO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AQ;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_BO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_BO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CLK;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_DO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A5Q;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_AMUX;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_AO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_AQ;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B5Q;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_BMUX;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_BO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_BO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_BQ;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_CLK;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_CO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_DO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_BO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_BO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CLK;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_DO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_CO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_DO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_AO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_AO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_AQ;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_BO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_BO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_CLK;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_CO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_CO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_DO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_DO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_AO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_AO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_BO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_CO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_CO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_DO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_DO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_AO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_AO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_BO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_BO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_BQ;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_CLK;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_CO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_DO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_DO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_AMUX;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_AO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_AO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_AQ;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_AX;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_BO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_BO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_CE;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_CLK;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_CO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_CO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_DO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_DO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_SR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_AO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_AO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_A_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_BO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_BO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_BQ;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_B_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_CLK;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_CO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_CO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_C_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_DO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_DO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X18Y116_D_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_AO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_AO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_A_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_BO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_BO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_B_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_CO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_CO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_C_XOR;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D1;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D2;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D3;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D4;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_DO5;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_DO6;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D_CY;
  wire [0:0] CLBLM_R_X13Y116_SLICE_X19Y116_D_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BMUX;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CLK;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_DO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_AO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_AO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_BO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_BO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_CO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_CO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_DO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_DO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_BO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_BO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CLK;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_DO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_DO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_AO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_AO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_BO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_BO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_CO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_CO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_DO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_DO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D_XOR;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_A;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_A1;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_A2;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_A3;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_A4;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_A5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_A6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_AO5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_AO6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_A_CY;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_A_XOR;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_B;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_B1;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_B2;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_B3;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_B4;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_B5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_B6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_BO5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_BO6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_B_CY;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_B_XOR;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_C;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_C1;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_C2;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_C3;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_C4;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_C5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_C6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_CO5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_CO6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_C_CY;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_C_XOR;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_D;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_D1;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_D2;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_D3;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_D4;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_D5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_D6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_DO5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_DO6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_D_CY;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X56Y115_D_XOR;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_A;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_A1;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_A2;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_A3;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_A4;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_A5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_A6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_AO5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_AO6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_A_CY;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_A_XOR;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_B;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_B1;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_B2;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_B3;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_B4;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_B5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_B6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_BO5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_BO6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_B_CY;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_B_XOR;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_C;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_C1;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_C2;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_C3;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_C4;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_C5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_C6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_CO5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_CO6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_C_CY;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_C_XOR;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_D;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_D1;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_D2;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_D3;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_D4;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_D5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_D6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_DO5;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_DO6;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_D_CY;
  wire [0:0] CLBLM_R_X37Y115_SLICE_X57Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AQ;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CLK;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CLK;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CLK;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CLK;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CLK;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CLK;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5Q;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CLK;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5Q;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CLK;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CLK;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CLK;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CLK;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5Q;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CLK;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CLK;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CLK;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CLK;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5Q;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CLK;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CLK;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CLK;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5Q;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CLK;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CLK;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CLK;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CLK;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CLK;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CLK;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5Q;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CLK;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CLK;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CLK;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CLK;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BMUX;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CLK;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CLK;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5Q;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A5Q;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A5Q;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AX;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CLK;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B5Q;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CLK;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CLK;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A5Q;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B5Q;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CLK;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AQ;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CLK;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CLK;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CLK;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CLK;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CLK;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CLK;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CLK;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CLK;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CLK;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CLK;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5Q;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CLK;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5Q;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5Q;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CLK;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CLK;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CLK;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5Q;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffdffffffdd)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_DLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffddfffdfffd)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddfffffffcffff)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_BLUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffcfffefffef)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000dccc0000cccc)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_ALUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_DQ),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_BQ),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfcddccf5f05500)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.I2(LIOB33_X0Y51_IOB_X0Y51_I),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000eac00000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I1(LIOB33_X0Y53_IOB_X0Y53_I),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_D5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f000f000f0)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_AO6),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f007777ffff)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_BO6),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h44cc44cc55ff55ff)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff44ff00000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_DQ),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_B5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffcfaaaa0a0a)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_DQ),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffce)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I3(CLBLL_L_X2Y114_SLICE_X1Y114_BO6),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.I5(CLBLL_L_X2Y113_SLICE_X1Y113_BO6),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00730050)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I4(LIOB33_X0Y67_IOB_X0Y68_I),
.I5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010001000110000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I4(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf050f050f050fcdc)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_DLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(LIOB33_X0Y67_IOB_X0Y67_I),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_BQ),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000320010)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeefffffffe)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_ALUT (
.I0(CLBLL_L_X2Y114_SLICE_X1Y114_DO6),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_CO6),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3ffffffcffffff)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000003300f3f0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I2(LIOB33_X0Y61_IOB_X0Y61_I),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000a000c)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00a00040)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbffffdfff)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044001010)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_DLUT (
.I0(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I3(LIOB33_X0Y55_IOB_X0Y55_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fff3ffff3f3f3f3)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffffffffffbf)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fff0000a040)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.Q(CLBLL_L_X4Y108_SLICE_X4Y108_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.Q(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.Q(CLBLL_L_X4Y108_SLICE_X4Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.Q(CLBLL_L_X4Y108_SLICE_X4Y108_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfffacccc0050)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_DQ),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_DQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2c0c0ffddffdd)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_BQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaeefb0000ccf3)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_BQ),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0b1a0ff000000)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_DO6),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.Q(CLBLL_L_X4Y108_SLICE_X5Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.Q(CLBLL_L_X4Y108_SLICE_X5Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.Q(CLBLL_L_X4Y108_SLICE_X5Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcf0f0fcfcf0f0f)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ff050ff4fc040c)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_DQ),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc000055aa)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_DO6),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc10fe32dc10dc10)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_AQ),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbfffffffff)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_D5Q),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200020002000a00)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_D5Q),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafaaaf888f888)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5550ccccfff0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_DO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00a0a00a0a)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(CLBLL_L_X2Y110_SLICE_X1Y110_AO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_DQ),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_CQ),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888f8f8800ffffff)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_C5Q),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_A5Q),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fe54fe54fe54)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003232ff00fafa)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbbbbbbbfbbbfbb)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_B5Q),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_DQ),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_BQ),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fa0aacacacac)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafaaaf888f888)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000c000c0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.Q(CLBLL_L_X4Y110_SLICE_X5Y110_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.Q(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.Q(CLBLL_L_X4Y110_SLICE_X5Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.Q(CLBLL_L_X4Y110_SLICE_X5Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h060a0a0a0a0a0a0a)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_A5Q),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_CQ),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_A5Q),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_DQ),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f09900cc00)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_CQ),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_AO6),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acfc0cfc0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8a8a8ffa8a8a8)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_BQ),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc008ccccc8c8c)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff030c0000030c)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_C5Q),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa8a8a8a8a8a8)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_BQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y110_SLICE_X16Y110_D5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfceefc00302230)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X13Y111_SLICE_X19Y111_BQ),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.Q(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.Q(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.Q(CLBLL_L_X4Y111_SLICE_X5Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.Q(CLBLL_L_X4Y111_SLICE_X5Y111_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aafcaafcaafc)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_BQ),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aafcaafcaafc)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_CQ),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff4400440044)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffa800fc00a8)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLL_L_X4Y110_SLICE_X5Y110_CQ),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88d8888888888888)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f404f404)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_CQ),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccccff00)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_CQ),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000c4c0c4c0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_CQ),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.Q(CLBLL_L_X4Y112_SLICE_X5Y112_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.Q(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.Q(CLBLL_L_X4Y112_SLICE_X5Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.Q(CLBLL_L_X4Y112_SLICE_X5Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300bbaabbaa)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8fcfc3030)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff008080ff000000)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_A5Q),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_A5Q),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_CQ),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_DQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacfcac0cfcfc0c0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.Q(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.Q(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000c0a0e0a0e)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3f330f00)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_BO6),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CQ),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff9fc0f0f090c)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_CQ),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300fcfc3030)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfefefcccceeee)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I3(1'b1),
.I4(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4fff4f4f44ff4444)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_CQ),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_BO6),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_AQ),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_CO6),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ccccf0f0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_CQ),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040404ff0404)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000033000a0a3b0a)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_CQ),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000800000)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_CO6),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d0cffff5d0c5d0c)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_DQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000400050000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_DQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_DO6),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeffeffffff)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0eeeeaaaa)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0aff0a0a)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(1'b1),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffdfffcfffc)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_CO6),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_A5Q),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdfffffffc)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_DO6),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_DO6),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_CO6),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7575ffff3030)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_DO6),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_DQ),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_DO6),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_BO6),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f444f44ffff4f44)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ff55fa50aa00)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_DQ),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_CQ),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffcfffcc)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_DO6),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_CO6),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff73ffffff50)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I2(LIOB33_X0Y65_IOB_X0Y66_I),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I4(CLBLM_R_X5Y117_SLICE_X6Y117_DO6),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_CQ),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff2ff00002222)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(LIOB33_X0Y65_IOB_X0Y65_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_A5Q),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbffeffffff)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3fff0fffbfffa)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_CQ),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I3(CLBLL_L_X4Y116_SLICE_X5Y116_CO6),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000800000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffafffbbffaa)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_A5Q),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfffcfffff3fff3)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_DO6),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000100)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.I1(CLBLL_L_X2Y113_SLICE_X1Y113_CO6),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffff40400000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdffffffffffeff)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfdfcf00005500)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafe)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010001000330010)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1100000011300030)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000004030003)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h002200220f2f0022)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_CLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffff33000000)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdefffefefffffff)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3ffc000f300c0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00de12cc00cc00)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_D5Q),
.I4(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.Q(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.Q(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.Q(CLBLM_L_X8Y106_SLICE_X10Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000fc0cfc0c)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_B5Q),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaaeeaa44004400)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y108_SLICE_X5Y108_BQ),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbabbba11101110)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.Q(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.Q(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.Q(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000010005000)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I4(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaaaea00500040)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hea40ea40ee44ee44)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_C5Q),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888888d8d8)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_CQ),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.Q(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.Q(CLBLM_L_X8Y107_SLICE_X11Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.Q(CLBLM_L_X8Y107_SLICE_X11Y107_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000af00af)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_DLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00a8000000a8)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_CQ),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff54ff5400540054)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_B5Q),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e1f0f000000044)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_ALUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.Q(CLBLM_L_X8Y108_SLICE_X10Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.Q(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.Q(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffe)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_DLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0f5a0e4a0e4)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_BQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc4ffc400c400c4)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_CQ),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafff0ccc0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_ALUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.Q(CLBLM_L_X8Y108_SLICE_X11Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.Q(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.Q(CLBLM_L_X8Y108_SLICE_X11Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.Q(CLBLM_L_X8Y108_SLICE_X11Y108_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaaafa00500050)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cacaff000a0a)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_CLUT (
.I0(CLBLM_L_X12Y112_SLICE_X17Y112_AQ),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_CQ),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fef0fe000e000e)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fe10fe10)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_AQ),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_CQ),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.Q(CLBLM_L_X8Y109_SLICE_X10Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.Q(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.Q(CLBLM_L_X8Y109_SLICE_X10Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333339fffff0ff)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00fef40e04)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffa800fc00a8)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_C5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fff0fff0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X11Y109_DO6),
.Q(CLBLM_L_X8Y109_SLICE_X11Y109_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.Q(CLBLM_L_X8Y109_SLICE_X11Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.Q(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.Q(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afac00330033)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_DLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y109_SLICE_X11Y109_A5Q),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0a0800000a08)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1a0b1a0e4a0e4)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.I2(CLBLM_L_X12Y112_SLICE_X17Y112_AQ),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00ff30fc)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_AQ),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.Q(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.Q(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.Q(CLBLM_L_X8Y110_SLICE_X10Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005555ffff5555)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heac0faf0faf0eac0)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CQ),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_DO6),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f60006f0f60006)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0055555050)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.Q(CLBLM_L_X8Y110_SLICE_X11Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.Q(CLBLM_L_X8Y110_SLICE_X11Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AQ),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_DO5),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cc00f0aaf0aa)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I2(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'habae0104aeae0404)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_BQ),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_AQ),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc55505550)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_CQ),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.Q(CLBLM_L_X8Y111_SLICE_X10Y111_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.Q(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff006c6cff00cccc)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cc00df00ec00)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I1(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_C5Q),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_CQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hea40ea40f5f5a0a0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.Q(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.Q(CLBLM_L_X8Y111_SLICE_X11Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.Q(CLBLM_L_X8Y111_SLICE_X11Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f000f0f87008)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc480c080c080c080)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4e4dd88dd88)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_BQ),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafff0ccc0)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_A5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_AQ),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_CQ),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeee00000eee0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_DQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafcfafc0a0c0a0c)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaefeae54045404)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_DQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y112_SLICE_X14Y112_BQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fefe5454)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.Q(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.Q(CLBLM_L_X8Y112_SLICE_X11Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00000eeee0000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01ba10ab01ba10)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_CQ),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_B5Q),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888dddd8888d8d8)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_C5Q),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5050cccc5050)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y113_SLICE_X17Y113_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0aaaaf0f0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5e4f5e4)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_BQ),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.I3(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00fcfcfc)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_DQ),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_CO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_DO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c5c0c0c5c5c0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff001414ff001414)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff6c0000006c)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fafac8c8)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_DQ),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_DO5),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_CO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_DO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f033aa00aacc)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_D5Q),
.I1(RIOB33_X105Y119_IOB_X1Y119_I),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f000aaf0aaff)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_DQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaf0f00a0a0000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_D5Q),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000200000002)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_ALUT (
.I0(RIOB33_X105Y119_IOB_X1Y119_I),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_BO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffc0cf000fc0c)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfff000f0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f6f688888888)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_DLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a3a0aca0aca0ac)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_DQ),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_DO5),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaccaaf0aacc)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_C5Q),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf005055555)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_BO5),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000008080000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_CLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_AO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888f5a0f5a0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I2(CLBLM_R_X11Y112_SLICE_X14Y112_DQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f30303f0f10001)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_A5Q),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_DO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa30aa33aa30)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_DLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_BQ),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f011444444)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_CLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_CQ),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afa0acacafa0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50aa00be14aa00)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_AO6),
.I5(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22000000cc00fc30)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_C5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0f000f00)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3faaffaaffaaff)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_B5Q),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_C5Q),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_AO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_BO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_CO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000ff00)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_CLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff4400440044)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fccf0cc00cc00)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_AO6),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0bf00000ff000000)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_D5Q),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_BO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_CO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_DO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0050505050)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afafafa0afac)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000a0aff00caca)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_BLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff004444ff00e4e4)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_ALUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_CLUT (
.I0(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_D5Q),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555545500000300)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff32ff1000320010)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d888d800f000f0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_B5Q),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_A5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.Q(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.Q(CLBLM_L_X10Y106_SLICE_X12Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.Q(CLBLM_L_X10Y106_SLICE_X12Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000eeee)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_CLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_CQ),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cd01cf03cd01)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_BLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff3000330030)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_CQ),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9009900990099009)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_DLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_A5Q),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_D5Q),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000011dd11dd)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_CLUT (
.I0(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_BQ),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000bbaa4455ffff)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.I2(1'b1),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_DQ),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff5ffffffff5ff5)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_ALUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_B5Q),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_DQ),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_CQ),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.Q(CLBLM_L_X10Y107_SLICE_X12Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_CQ),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000a4e00005f1b)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_CQ),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_DQ),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f06050605)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_BQ),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_AQ),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_D5Q),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfdccfd00310031)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.Q(CLBLM_L_X10Y107_SLICE_X13Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.Q(CLBLM_L_X10Y107_SLICE_X13Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c553c3c3caa)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_DLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_A5Q),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_CQ),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_CO5),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000055445544)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_CQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffc00fc)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_BQ),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_DQ),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc9cc00aa00aa)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_ALUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.Q(CLBLM_L_X10Y108_SLICE_X12Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.Q(CLBLM_L_X10Y108_SLICE_X12Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.Q(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f050f050f0d0f0d)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_DLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cc00aaaa)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_CLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0ccfffff088)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_BQ),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00dc1033333030)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_ALUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.Q(CLBLM_L_X10Y108_SLICE_X13Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5affffffff5a5a)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_DLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_CQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_A5Q),
.I5(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699669999669966)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_CLUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_BQ),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_CQ),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4040101004040101)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_BLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb888bbbbb8888888)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_CQ),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.Q(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000a0a)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ccfcaaaaaaaa)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_CLUT (
.I0(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_CQ),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb00ff5500000000)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffc00fc)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.Q(CLBLM_L_X10Y109_SLICE_X13Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.Q(CLBLM_L_X10Y109_SLICE_X13Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ccffffffff33cc)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y109_SLICE_X18Y109_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_CQ),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0900000900000000)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_CLUT (
.I0(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_A5Q),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afafacac)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_BLUT (
.I0(CLBLM_R_X13Y109_SLICE_X18Y109_CQ),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf000aaaafc00)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_ALUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_A5Q),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_CQ),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.Q(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.Q(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.Q(CLBLM_L_X10Y110_SLICE_X12Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00e0e0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_DQ),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc00fc00fc00)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_CLUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_BQ),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0b1b1e4e4)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_BQ),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.I3(1'b1),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dc10dd11dc10)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88d888888888)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_AQ),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef45af05ea40aa00)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_CQ),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X13Y109_SLICE_X18Y109_BQ),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eeeef0f04444)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_DQ),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa30aa33aa30)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_ALUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X12Y111_DO5),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccff005050)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_CQ),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11cc00dd11cc00)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_AQ),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaa00c0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_DQ),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_BQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ffaaaa00f0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_DO5),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b88888ffcc3300)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccaaf0aa00)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_A5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y115_SLICE_X14Y115_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888d8d8a0a0f5a0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_CQ),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_BQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000fa00fa)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.Q(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccfcfdddddfdf)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_DLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffa0e4a0e4)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050505540404055)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_BLUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_DQ),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafff0ffaaffc0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_ALUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.Q(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.Q(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.Q(CLBLM_L_X10Y112_SLICE_X13Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffccaaaaf0c0)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_DQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafe0054fefe5454)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_DQ),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a0a0ffcc0000)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_DQ),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_BQ),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddd8888888d8)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_DQ),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X11Y112_SLICE_X14Y112_BQ),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0a0a0f0c0f0c)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_DLUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_DQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_AQ),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00dd11dd11cc00)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hba10ba10ba10ba10)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_DQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc55cc50cc50)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_A5Q),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_AO6),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfffffffcff)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000020)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_CQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cacac0c0c5c5)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_BLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_BO5),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffccc3000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_DO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8bbbbb8b88888)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_DLUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_DQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5e4a0a0f5e4)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_CQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_DQ),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_CQ),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafcfafcfafcfaf0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefeeedcdcdccc)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_A5Q),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_CO5),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_AO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff12ff1200120012)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_DLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_CO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00acacacac)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_CLUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hababaeae01010404)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_CQ),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfecccc00320000)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_ALUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_CO5),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_DO5),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_BO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_CO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_DO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0aaccaacc)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_DLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_C5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0f0f000aa)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_C5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_D5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbffff0f0b0f0f)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y118_SLICE_X11Y118_BO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdffff0f0d0f0f)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y118_SLICE_X11Y118_BO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X13Y115_AO6),
.Q(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.Q(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.Q(CLBLM_L_X10Y115_SLICE_X13Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_DLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_CQ),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_DQ),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_DQ),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe5554ffaa5500)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_BO6),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe5554aaae0004)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X12Y114_SLICE_X17Y114_CQ),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_DQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccccfcecfcec)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_CO5),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_AO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_CO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0ffffaa00)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404cfcfc0c0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_BQ),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0aca00000aca)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_BLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbbbbb8bbbb)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_L_X8Y118_SLICE_X11Y118_BO6),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_AO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aaaa56665666)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_CQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00fa00ff00ea0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_BLUT (
.I0(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_CQ),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccceeddc00022110)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f044444444)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000fc0cfc0c)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y116_SLICE_X18Y116_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f07722f0f05500)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_BLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_CQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff007575ff002020)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_ALUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555777f5555777f)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_DLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_CQ),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300ffff0100ffff)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_D5Q),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_CO6),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_CQ),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeee0a000a00)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_D5Q),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e2e2ff00f3f3)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_BO5),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_CO5),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0fff00f00)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_CLUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y143_IOB_X1Y144_I),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00ccf0f0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_BLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1f5a0e4b1b1a0a0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_C5Q),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa55a9aaaa5555)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_DLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff1b0000ffff)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa000000005050)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I3(1'b1),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h444544450000fffe)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_D5Q),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.R(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.R(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55fd55ff55ff)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_DLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_D5Q),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033133212)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_D5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100001000)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf30051ff5d550cbb)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_D5Q),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_BO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d0d0f0f0c0f0f0f)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_DLUT (
.I0(CLBLM_L_X12Y118_SLICE_X16Y118_AO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I3(CLBLM_L_X12Y118_SLICE_X16Y118_AO5),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000003030)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_L_X12Y118_SLICE_X16Y118_AO5),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffc600c6)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_BLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f008f8f4f004f4f)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2c3d2c3d2c3d2c3)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f300f3f3f300f3)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I5(CLBLM_L_X10Y120_SLICE_X13Y120_CO6),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0eef0aaf0ee)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_ALUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333ffaa5500)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_A5Q),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000f3f3f3f3)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfffc30303330)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777fffff0000000)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_ALUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_C5Q),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_B5Q),
.I2(RIOB33_X105Y139_IOB_X1Y140_I),
.I3(RIOB33_X105Y141_IOB_X1Y141_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.Q(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y107_SLICE_X16Y107_BO6),
.Q(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y107_SLICE_X16Y107_CO6),
.Q(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hecccccccecccffff)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaafe00540054)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y111_SLICE_X19Y111_AQ),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f808f404)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_BLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac0c0aaaaff00)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_ALUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.Q(CLBLM_L_X12Y108_SLICE_X16Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.Q(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a05050a050a0a05)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_DLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00010c0d03020f0e)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_CLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_BO5),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_A5Q),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdd3311fcdc3010)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_BLUT (
.I0(CLBLM_L_X12Y108_SLICE_X16Y108_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I4(CLBLM_R_X11Y113_SLICE_X15Y113_DQ),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa33aa30aa30)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_ALUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_A5Q),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y108_SLICE_X17Y108_AO6),
.Q(CLBLM_L_X12Y108_SLICE_X17Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y108_SLICE_X17Y108_BO6),
.Q(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffaaffaa)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_DLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y112_SLICE_X17Y112_AQ),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_CLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y108_SLICE_X11Y108_CQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y109_SLICE_X18Y109_BQ),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff0ffc0c)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_AQ),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd500d5ff800080)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y108_SLICE_X17Y108_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_AQ),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y109_SLICE_X16Y109_AO6),
.Q(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6fffff6f6fffff6)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_DLUT (
.I0(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_CQ),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_CLUT (
.I0(CLBLM_L_X12Y108_SLICE_X17Y108_AQ),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_CQ),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I3(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_CQ),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc0002fffd)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_BLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I4(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0041410000)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_DO5),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0000fbff0000fb)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_DLUT (
.I0(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_CO6),
.I2(CLBLM_L_X12Y108_SLICE_X17Y108_DO6),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.I4(CLBLM_R_X13Y109_SLICE_X18Y109_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44eeeeee444444)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_CLUT (
.I0(CLBLM_L_X12Y111_SLICE_X17Y111_CO5),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.I4(CLBLM_R_X13Y109_SLICE_X18Y109_AQ),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_BO6),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffef)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_BLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I1(CLBLM_L_X12Y112_SLICE_X17Y112_AQ),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_CO6),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_AQ),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0d00000f0e00000)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_ALUT (
.I0(CLBLM_L_X12Y109_SLICE_X17Y109_DO6),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_DO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_R_X11Y109_SLICE_X15Y109_CO6),
.I4(CLBLM_L_X12Y111_SLICE_X17Y111_CO5),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.Q(CLBLM_L_X12Y110_SLICE_X16Y110_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X16Y110_AO6),
.Q(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.Q(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X16Y110_CO6),
.Q(CLBLM_L_X12Y110_SLICE_X16Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X16Y110_DO6),
.Q(CLBLM_L_X12Y110_SLICE_X16Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaacccc)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_DLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_AQ),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_D5Q),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cacaff000a0a)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_CLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_CQ),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd500d5ff800080)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_CQ),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdddeccc31112000)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_AQ),
.I5(CLBLM_L_X12Y114_SLICE_X16Y114_CQ),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X17Y110_AO6),
.Q(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X17Y110_BO6),
.Q(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X17Y110_CO6),
.Q(CLBLM_L_X12Y110_SLICE_X17Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0faf0fef0fef0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_BO5),
.I2(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afa0a0a0aca0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_CLUT (
.I0(CLBLM_R_X13Y109_SLICE_X18Y109_AQ),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_AQ),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d580d580)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300fedc3210)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_CQ),
.I4(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y111_SLICE_X16Y111_BO5),
.Q(CLBLM_L_X12Y111_SLICE_X16Y111_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y111_SLICE_X16Y111_AO6),
.Q(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y111_SLICE_X16Y111_BO6),
.Q(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaa5a5aaaaa5a5)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_DLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I3(1'b1),
.I4(CLBLM_L_X12Y113_SLICE_X16Y113_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_DO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffafffffffa)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_CLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I4(CLBLM_R_X13Y112_SLICE_X18Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_CO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaacccc)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_BLUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I1(CLBLM_R_X11Y116_SLICE_X15Y116_CQ),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_BO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff12ff2400120024)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_ALUT (
.I0(CLBLM_L_X12Y111_SLICE_X16Y111_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_C5Q),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_AO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y111_SLICE_X17Y111_AO6),
.Q(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y111_SLICE_X17Y111_BO6),
.Q(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffccffcc)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_BO5),
.I4(1'b1),
.I5(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_DO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f0f0f088000000)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_CLUT (
.I0(CLBLM_R_X13Y111_SLICE_X19Y111_AQ),
.I1(CLBLM_R_X13Y111_SLICE_X19Y111_BQ),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_BQ),
.I4(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_CO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecececfca0a0a0f0)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_BLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y118_SLICE_X16Y118_BO6),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I5(CLBLM_R_X13Y115_SLICE_X18Y115_BQ),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_BO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3000aaaa0300)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_ALUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_CQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I2(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y111_SLICE_X17Y111_CO6),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_AO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X15Y112_BO6),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X16Y112_CO6),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X16Y112_AO6),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X16Y112_BO6),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa000004444)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_DLUT (
.I0(CLBLM_L_X12Y112_SLICE_X17Y112_BQ),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y112_SLICE_X16Y112_A5Q),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_DO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacafafac0000ff00)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_CLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_CO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f40104f0f40004)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I1(CLBLM_L_X12Y112_SLICE_X16Y112_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y112_SLICE_X16Y112_DO5),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_CQ),
.I5(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_BO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31ec20dd11cc00)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_AO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X17Y112_AO6),
.Q(CLBLM_L_X12Y112_SLICE_X17Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X17Y112_BO6),
.Q(CLBLM_L_X12Y112_SLICE_X17Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X17Y112_CO6),
.Q(CLBLM_L_X12Y112_SLICE_X17Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0a0a0f0c0f0c)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_DLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_DQ),
.I1(CLBLM_L_X12Y112_SLICE_X17Y112_CQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I3(CLBLM_R_X13Y109_SLICE_X18Y109_DQ),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_DO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afa0a0a0aca0)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.I1(CLBLM_L_X12Y112_SLICE_X17Y112_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_CO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aabe0014)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y112_SLICE_X17Y112_BQ),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_CO5),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I5(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_BO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5cca0cc55cc00)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I1(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.I2(CLBLM_L_X12Y112_SLICE_X17Y112_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y110_SLICE_X16Y110_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_AO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X16Y113_AO6),
.Q(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X16Y113_BO6),
.Q(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X16Y113_CO6),
.Q(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X16Y113_DO6),
.Q(CLBLM_L_X12Y113_SLICE_X16Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa00aa0faa00)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_DLUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_DO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaffaa40405500)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I5(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_CO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00fc0c)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_DQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_BO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccffccf0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_BQ),
.I2(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_AO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X17Y113_AO6),
.Q(CLBLM_L_X12Y113_SLICE_X17Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X17Y113_BO6),
.Q(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X17Y113_CO6),
.Q(CLBLM_L_X12Y113_SLICE_X17Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_DO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffacacffffaca0)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_CLUT (
.I0(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.I1(CLBLM_L_X12Y113_SLICE_X17Y113_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_CO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecec2020ecec2020)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y112_SLICE_X18Y112_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_BO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0fff066)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_ALUT (
.I0(CLBLM_L_X12Y113_SLICE_X17Y113_AQ),
.I1(CLBLM_L_X12Y115_SLICE_X17Y115_BO6),
.I2(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.I5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_AO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X16Y114_AO6),
.Q(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X16Y114_BO6),
.Q(CLBLM_L_X12Y114_SLICE_X16Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.Q(CLBLM_L_X12Y114_SLICE_X16Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X16Y114_DO6),
.Q(CLBLM_L_X12Y114_SLICE_X16Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fc30ee22ee22)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_DLUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_DQ),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_DQ),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I5(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_DO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ee44fa50fa50)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_CQ),
.I2(CLBLM_R_X13Y116_SLICE_X18Y116_BQ),
.I3(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I5(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_CO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0074743030)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I1(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_CQ),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.I4(CLBLM_L_X12Y114_SLICE_X16Y114_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_BO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0e2e2e2e2)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_AO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X17Y114_AO6),
.Q(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X17Y114_BO6),
.Q(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X17Y114_CO6),
.Q(CLBLM_L_X12Y114_SLICE_X17Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haafbffaeaaffffaa)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_DLUT (
.I0(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.I1(CLBLM_R_X13Y115_SLICE_X18Y115_CO6),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I3(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.I4(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I5(CLBLM_L_X12Y114_SLICE_X16Y114_BQ),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_DO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ccf0aaf0aa)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_CLUT (
.I0(CLBLM_R_X13Y114_SLICE_X18Y114_AQ),
.I1(CLBLM_L_X12Y114_SLICE_X17Y114_CQ),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I5(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_CO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5f5e4e4)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y115_SLICE_X17Y115_AO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_BQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.I5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_BO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0aaf0aa)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_ALUT (
.I0(CLBLM_L_X12Y114_SLICE_X17Y114_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_AO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y110_SLICE_X16Y110_DQ),
.Q(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.R(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_DLUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I2(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I3(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_BO5),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_CLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_CO5),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.I4(CLBLM_R_X13Y115_SLICE_X19Y115_AO6),
.I5(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333233133333333)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_BLUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_BO5),
.I1(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I5(CLBLM_L_X12Y114_SLICE_X16Y114_CQ),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h444544450000fffe)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I1(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_CO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff0fef0fff)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_DLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffffffffffffff)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_CLUT (
.I0(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I1(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_BO5),
.I3(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I4(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff02ff0aff02)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_BLUT (
.I0(CLBLM_R_X13Y114_SLICE_X18Y114_AQ),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_DO6),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I3(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.I4(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.I5(CLBLM_L_X12Y115_SLICE_X17Y115_CO6),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h54ab55aa50af55aa)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_ALUT (
.I0(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_DO6),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I3(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.I5(CLBLM_L_X12Y115_SLICE_X17Y115_CO6),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X16Y116_AO6),
.Q(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3fcf6fcf6)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_DLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_BQ),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I2(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_DO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0057ffff03030303)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(CLBLM_R_X13Y115_SLICE_X19Y115_AO6),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_CO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h85a5c5f5aaaaa0a0)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_BO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000030123012)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_CO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_BO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_AO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X17Y116_AO6),
.Q(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X17Y116_BO6),
.Q(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4455bbaa4555baaa)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_DLUT (
.I0(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I2(CLBLM_R_X13Y117_SLICE_X18Y117_CO6),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I5(CLBLM_L_X12Y118_SLICE_X17Y118_BO6),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_DO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222330022223300)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_CLUT (
.I0(CLBLM_L_X12Y118_SLICE_X17Y118_BO6),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y117_SLICE_X18Y117_CO6),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_CO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f404f505f101)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_BLUT (
.I0(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I4(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.I5(CLBLM_L_X12Y117_SLICE_X17Y117_CO6),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_BO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffee00ee)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_DO6),
.I1(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_AO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_AO6),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0d08f8f7070af8c)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_DLUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_CO5),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_CO6),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_DO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00200000ffddffff)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_CLUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I1(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_CO6),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_CO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300020000)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_BLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.I1(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I2(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_BO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1c0d1c0d1c0d1c0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_ALUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_AO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X17Y117_AO6),
.Q(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008080808080)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_DLUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I2(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_DO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0b0e0f0f0f0f0f)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_CLUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I1(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I2(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.I3(CLBLM_R_X13Y117_SLICE_X18Y117_DO6),
.I4(CLBLM_L_X12Y117_SLICE_X17Y117_DO6),
.I5(CLBLM_L_X12Y114_SLICE_X16Y114_DQ),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_CO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a4b5a5a5a1e5a5a)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_BLUT (
.I0(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I4(CLBLM_R_X13Y116_SLICE_X18Y116_BQ),
.I5(CLBLM_L_X12Y116_SLICE_X16Y116_BO5),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_BO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000fffc3330)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.I3(CLBLM_L_X12Y117_SLICE_X17Y117_BO6),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_AQ),
.I5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_AO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_DO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_CO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303033333333)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_BO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000004)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_ALUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I4(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_AO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.Q(CLBLM_L_X12Y118_SLICE_X17Y118_AQ),
.R(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001100)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_DLUT (
.I0(CLBLM_L_X12Y113_SLICE_X17Y113_AQ),
.I1(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y117_SLICE_X18Y117_DO6),
.I4(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_DO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ffffffffffffff)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_CLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I1(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.I4(CLBLM_L_X12Y117_SLICE_X17Y117_DO6),
.I5(CLBLM_L_X12Y113_SLICE_X17Y113_AQ),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_CO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X17Y117_DO6),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I2(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.I3(CLBLM_L_X12Y113_SLICE_X17Y113_AQ),
.I4(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.I5(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_BO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fff70800fff30c)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_ALUT (
.I0(CLBLM_L_X12Y118_SLICE_X17Y118_DO6),
.I1(CLBLM_L_X12Y114_SLICE_X17Y114_CQ),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I3(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.I4(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.I5(CLBLM_L_X12Y118_SLICE_X17Y118_CO6),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_AO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0caa0caaaaffff)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_ALUT (
.I0(CLBLM_L_X12Y118_SLICE_X17Y118_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.Q(CLBLM_R_X3Y108_SLICE_X2Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y108_SLICE_X2Y108_BO6),
.Q(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff80ff80008000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_AQ),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_BQ),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00004000ffffb3ff)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_CLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_AQ),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_BQ),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f0f1f004000100)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5005cccc0000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_BQ),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_AQ),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.Q(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333ffffffff)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff77770fff0000)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_CLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fffffff)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_BLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_AQ),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_BQ),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff444000004440)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_DQ),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_BO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fffffff)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfef000000aa00aa)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_D5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cc330000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I3(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff008080c4c4)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_DO6),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.Q(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X3Y109_BO6),
.Q(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.Q(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff33ffffff)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacaca3aca0a0a0a0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_BQ),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heafa4050baaa1000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I4(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000030b830b8)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.Q(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.Q(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c000003333ffff)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cf03cc00ce02)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00dd11dc10)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.Q(CLBLM_R_X3Y110_SLICE_X3Y110_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.Q(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.Q(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.Q(CLBLM_R_X3Y110_SLICE_X3Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.Q(CLBLM_R_X3Y110_SLICE_X3Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff0033d1d1d1d1)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_BQ),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888b8b8b8b8)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff3300000033)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_C5Q),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_DQ),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffa0aaaaa0a0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.Q(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.Q(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb1111aaaa0000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_CQ),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hea00aa00c0000000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.Q(CLBLM_R_X3Y111_SLICE_X3Y111_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.Q(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.Q(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.Q(CLBLM_R_X3Y111_SLICE_X3Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaff77ff77)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000f505f000)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ee44fa50ee44)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_CQ),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fa50ba10fa50)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_BQ),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.Q(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccff595aa6a5)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0bbb0bbb3cc3c33c)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaa69966996)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff030003ff300030)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00cfccafaaefee)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd00cf00dd00ff00)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I3(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030cccc0000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y111_SLICE_X12Y111_CQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffc300000fc30)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_A5Q),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0022002200ff0022)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I2(1'b1),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8ffa8a8a8a8a8)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_CQ),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000eeee)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3ffaaaac000)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h003b003b000a000a)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I2(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3030baba)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010111000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_DQ),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafbfafaf00330000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_DQ),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff33f3ffff00f0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff2f22)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I5(CLBLL_L_X2Y114_SLICE_X1Y114_DO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h040404040404ff04)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccaaffaa00)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeeffffffff)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_DO6),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff2f2fffff2222)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000008c00af)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_BO6),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50dc50dcffff50dc)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_CO6),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffffffffffdf)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e4e4ff00e4e4)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8ddddd8d88888)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fefe00005454)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_BQ),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0c000c)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff50ffffffdc)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I2(LIOB33_X0Y63_IOB_X0Y63_I),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_BO6),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_DO6),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefffffffefffeff)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_DO6),
.I2(CLBLL_L_X2Y114_SLICE_X1Y114_AO6),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000008000000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_CLUT (
.I0(LIOB33_X0Y71_IOB_X0Y71_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffeefe)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_BLUT (
.I0(CLBLL_L_X2Y117_SLICE_X1Y117_DO6),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_DO6),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfdfcfcf00550000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_C5Q),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000abaa0300)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I5(CLBLL_L_X2Y117_SLICE_X1Y117_CO6),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000d000e000d00)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faf0fafcfefcfe)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_DLUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I3(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000030ba30ba)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_CLUT (
.I0(LIOB33_X0Y69_IOB_X0Y70_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020003000200000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y57_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaf0fffffefc)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I4(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I5(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefffef)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_DLUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_CLUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.I5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff7f)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_BLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.I3(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'habaaaababaaaaaaa)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000c555d000c)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.I4(LIOB33_X0Y59_IOB_X0Y59_I),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000050735050)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(LIOB33_X0Y53_IOB_X0Y54_I),
.I3(CLBLL_L_X2Y117_SLICE_X1Y117_CO6),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000000000000)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000080000)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000101f101)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1c0c0c0c0c0c0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffff00400004)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffffeffffff)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7f7ffffffbfb)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(1'b1),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X8Y107_CO5),
.Q(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.Q(CLBLM_R_X5Y107_SLICE_X7Y107_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.Q(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.Q(CLBLM_R_X5Y107_SLICE_X7Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.Q(CLBLM_R_X5Y107_SLICE_X7Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X7Y107_DO6),
.Q(CLBLM_R_X5Y107_SLICE_X7Y107_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000afa0afa0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_A5Q),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fcf0fc000c000c)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_D5Q),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cf000fc0c)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aafcaa30)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_ALUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_BQ),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.Q(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.Q(CLBLM_R_X5Y108_SLICE_X6Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.Q(CLBLM_R_X5Y108_SLICE_X6Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.Q(CLBLM_R_X5Y108_SLICE_X6Y108_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31ff33ec20cc00)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_DQ),
.I3(CLBLM_R_X13Y109_SLICE_X18Y109_BQ),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a0f5f5a0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_BQ),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_BQ),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00a8000000a8)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_BLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_BQ),
.I2(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_A5Q),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a0a0ff00f0f0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.Q(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.Q(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000545400005555)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_CLUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fcfccccc)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f30003f3f00300)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00fe54fe54)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f5f5e4e4a0a0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_C5Q),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f00500f4f00400)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y108_SLICE_X14Y108_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8a8a8ffa8a8a8)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.Q(CLBLM_R_X5Y109_SLICE_X7Y109_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.Q(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffffffffffffff)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_DQ),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_BQ),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000dffffffff)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_A5Q),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_A5Q),
.I3(LIOB33_X0Y53_IOB_X0Y53_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0af808aaaa8888)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X13Y109_SLICE_X18Y109_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_AQ),
.I4(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4a0e4e4f5b1f5f5)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_A5Q),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.I5(LIOB33_X0Y53_IOB_X0Y53_I),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.Q(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.Q(CLBLM_R_X5Y110_SLICE_X6Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000000)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_BQ),
.I5(CLBLL_L_X4Y108_SLICE_X5Y108_BQ),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffaf00f000f0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0033aaaa00cc)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaafa0000aafa)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.Q(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_DO6),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffdfffff)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_DQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_BQ),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00f0f0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffffff)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_CQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_BQ),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00aa00aa00)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffee440000ee44)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_AQ),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff007575ff003030)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.Q(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.Q(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.Q(CLBLM_R_X5Y111_SLICE_X7Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa00030000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haeeefeee04445444)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0c0c0cfc0c0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f202f101f202)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.Q(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.Q(CLBLM_R_X5Y112_SLICE_X6Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_CQ),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_BQ),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_CQ),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa00fa00ff00cc00)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_DQ),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f3f000030300)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c5c5c0c0caca)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_CQ),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.Q(CLBLM_R_X5Y112_SLICE_X7Y112_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.Q(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_A5Q),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_C5Q),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.I3(CLBLM_R_X5Y119_SLICE_X6Y119_A5Q),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_C5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_C5Q),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeefffffffe)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_A5Q),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_A5Q),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fa0afa0a)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50dc50dc50dc50dc)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_CQ),
.I3(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000500040000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_DQ),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff005454fcfc)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaeffaa04045500)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_CO6),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f55dfdd0f00cfcc)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f055fff0f044cc)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeafaeaf0c0f0c0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_DQ),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc0000fff0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_BQ),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0aff0aff0a)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_DLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_C5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000c0a)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_CLUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafaca0a0a0a0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_C5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe2ffaa00e200aa)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_B5Q),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I5(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_BO6),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3f3f3f3f3)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0affff0a0a0a0a)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44f5f5a0a0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_A5Q),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0003030c0c)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_DQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000faf000000aa)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff4f44)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_BQ),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_AQ),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff03ff00ff0bff0a)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(LIOB33_X0Y65_IOB_X0Y66_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_BO6),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.I5(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeffffeffff)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.Q(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X7Y115_BO6),
.Q(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff75ff30ff75ff30)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a02000008000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_CQ),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_DO6),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f00800f0f00000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_DQ),
.I5(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0aff0ffa0af000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_DQ),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000ccaa)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0bb88bb88)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_AQ),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbfffffffff7)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0e4a0f5a0e4)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffcccccc)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f5ccccf0a0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_A5Q),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaafa222222f2)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005522ffffffbb)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f03030ffffff33)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ccccfafa)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_A5Q),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_A5Q),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X7Y117_AO5),
.Q(CLBLM_R_X5Y117_SLICE_X7Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X7Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdfff)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_DLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff3bff0a)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_BO6),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000000000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaf0f0ff00)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_ALUT (
.I0(RIOB33_X105Y127_IOB_X1Y127_I),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffeffffffff)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(1'b1),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000000000000)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5fffa000)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I4(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaafaaa3c00f000)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_ALUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_BO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_CO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_DLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_A5Q),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe3caa00eeccaa00)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_A5Q),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000014001400)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_BLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff004848)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_CLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_A5Q),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff00080808080)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_CO6),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888b888888b888)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_CO6),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.Q(CLBLM_R_X7Y106_SLICE_X8Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.Q(CLBLM_R_X7Y106_SLICE_X8Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.Q(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.Q(CLBLM_R_X7Y106_SLICE_X8Y106_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888ddd88888)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_AQ),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_DQ),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaeafae05040504)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5a0e4a0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_BQ),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffb0b00000b0b0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_CQ),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X9Y106_BO5),
.Q(CLBLM_R_X7Y106_SLICE_X9Y106_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.Q(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.Q(CLBLM_R_X7Y106_SLICE_X9Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X9Y106_CO6),
.Q(CLBLM_R_X7Y106_SLICE_X9Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000003003fccf)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_B5Q),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef45ea40ee44ee44)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_CQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444fa50fa50)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_B5Q),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c0c5c5c5c0c5)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_DO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.Q(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.Q(CLBLM_R_X7Y107_SLICE_X8Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000110011)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_DLUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BQ),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h10101010afaa0500)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54fe54aa00)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_BQ),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb33ba30aa00aa00)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_DO5),
.I5(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.Q(CLBLM_R_X7Y107_SLICE_X9Y107_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.Q(CLBLM_R_X7Y107_SLICE_X9Y107_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.Q(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.Q(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffeeee)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_C5Q),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaa200005555)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ee44ee44)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaa0000)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_ALUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.Q(CLBLM_R_X7Y108_SLICE_X8Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.Q(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee2233333f3f)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_DLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_DQ),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a3a3acac)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_CLUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc00fc00fc00)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_BQ),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00ccccfa50)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_AQ),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0b0f0f0b0b0f0a0)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_DLUT (
.I0(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I4(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000efafaaaa)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_CLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_DQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000faf80000f2f0)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_AQ),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_DQ),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000ffffffefe)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_ALUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I2(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.Q(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.Q(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e0e0e0e0e0c5e0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5577557757725577)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_DQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404f000f000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_DQ),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aac0aaffaacc)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_A5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.Q(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.Q(CLBLM_R_X7Y109_SLICE_X9Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa55555aaa55555)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc900c9ffc900c9)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_DO5),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_CQ),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'habab0101baba1010)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hba10ab01ba10ab01)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_AQ),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.Q(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0f00ff00f0ff0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_DQ),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0010ffff0010)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0069960000699600)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff600060ff600060)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(CLBLM_R_X7Y108_SLICE_X9Y108_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.Q(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.Q(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffefffefff)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444cc4c44440000)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f000f044f000)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_DQ),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaafcaa00)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_A5Q),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_BQ),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.Q(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.Q(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.Q(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f1fffff0f0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_CO6),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_B5Q),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00de12de12)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000c3c3)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccff0f0f)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_DQ),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_B5Q),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.Q(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0e)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_BQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_DQ),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_B5Q),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc5cfc0c0cac0)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c6996c3cc996633)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_CQ),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_DO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_DQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc0f0cfaf80a08)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_BQ),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.Q(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.Q(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffbfb)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_C5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_C5Q),
.I3(1'b1),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_B5Q),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff888d0000f0f0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffcc00cc)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafff000f0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaa00cc00cc)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_C5Q),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h010000000e0f0f0f)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_C5Q),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_B5Q),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffef0000cfcf)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_D5Q),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11aa00ba10aa00)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_DQ),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(CLBLM_R_X11Y112_SLICE_X14Y112_DQ),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50ee44ee44)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_DQ),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fcaaaafcfc)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddddddd8888888)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_DQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefeeedcdcdccc)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_C5Q),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc55cc55cc00)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_BQ),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccfa00fa00)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I2(CLBLM_L_X10Y111_SLICE_X12Y111_D5Q),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0ccf0cc)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_CQ),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00cccc5050)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_DQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1c0d1c0fcfc3030)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fc30303030)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e4e4cccc)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.Q(CLBLM_R_X7Y114_SLICE_X9Y114_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.Q(CLBLM_R_X7Y114_SLICE_X9Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.Q(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X9Y114_CO6),
.Q(CLBLM_R_X7Y114_SLICE_X9Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000808000008000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044ccffcc00)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_CQ),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa03aa0faa0caa00)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(CLBLM_L_X12Y111_SLICE_X16Y111_B5Q),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000055505550)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I1(1'b1),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_CQ),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_AQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_BO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_CO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000c800000008)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_DO6),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0eca0eca0eca0ec)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_DQ),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf0fff000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_BQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffaaaaaa)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_BO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_CO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff20ff2000200020)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_DQ),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fefe5454)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000fcfc)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafafafacaf)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_B5Q),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff004444ccccf0f0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaa3c00eeaacc00)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaa0f00faaaf000)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff115533ff)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55550000f7d5f3c0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_CLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_L_X12Y111_SLICE_X16Y111_B5Q),
.I3(CLBLM_R_X13Y115_SLICE_X18Y115_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h575f77ffc0000000)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff33fc30)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_DO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_CO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaac000c000)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_DLUT (
.I0(RIOB33_X105Y127_IOB_X1Y127_I),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaa3300eeaacc00)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaa3c00eeaacc00)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0c0c0cffc0c0c0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_DO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee5044faee5044)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_A5Q),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I4(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3a0b3a055550000)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffcc00cc)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0ffc0cfc0c)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_C5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_BO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_CO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_DLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_AQ),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccaaccaa)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_B5Q),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f6f0f000060000)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_A5Q),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_A5Q),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fc30fc30)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005500000000)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000050f5f5f5f5)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(1'b1),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00afafff00fafa)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0000000000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00dc1010101010)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_BLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc00cc50cc00)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_ALUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0ccccccf0f0)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_D5Q),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_DO5),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d00000dfff2f2ff)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_B5Q),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_BLUT (
.I0(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00f0fe4b14e1b)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_ALUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc5a5a)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_DLUT (
.I0(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_A5Q),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_CO5),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcffffaa9aaaaa)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbff0400ff33ff33)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_BLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa9aaa00000f0f)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_ALUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_BQ),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.Q(CLBLM_R_X11Y107_SLICE_X15Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.Q(CLBLM_R_X11Y107_SLICE_X15Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3faaaa9aaa)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_DLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_BQ),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00008800f0b4f0f0)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_CLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_A5Q),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888b8b8b8b8)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_BLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22cc00cc00)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_ALUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_DQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.Q(CLBLM_R_X11Y108_SLICE_X14Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f550f99)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_DLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_AQ),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000335a3355)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_CLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_A5Q),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_AQ),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaa6ffffff0f)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ccccf0ff)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_AQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.Q(CLBLM_R_X11Y108_SLICE_X15Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_DLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_CQ),
.I1(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cc3c3c3c33c3c)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AQ),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_AQ),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_AQ),
.I3(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11bb11ba10ba10)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_AQ),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_CQ),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.Q(CLBLM_R_X11Y109_SLICE_X14Y109_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.Q(CLBLM_R_X11Y109_SLICE_X14Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.Q(CLBLM_R_X11Y109_SLICE_X14Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f5500000f66)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_DQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_DQ),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00dc10cc00)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I4(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb88b800000f0f)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccffcc0f)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_DO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ddbbee77ddbbee)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_DLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_AQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y112_SLICE_X17Y112_AQ),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff3c3c)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y109_SLICE_X15Y109_DO6),
.I5(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0fcfc)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_DQ),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_BQ),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_BQ),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_BO5),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00facccc00fa)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_DLUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_AQ),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_A5Q),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_DQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11aa00bb11aa00)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f00aaaa0c00)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_BLUT (
.I0(CLBLM_L_X12Y113_SLICE_X17Y113_CQ),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_AQ),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222f3c0f3c0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_A5Q),
.I4(CLBLM_R_X11Y110_SLICE_X15Y110_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.Q(CLBLM_R_X11Y110_SLICE_X15Y110_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.Q(CLBLM_R_X11Y110_SLICE_X15Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X15Y110_BO6),
.Q(CLBLM_R_X11Y110_SLICE_X15Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.Q(CLBLM_R_X11Y110_SLICE_X15Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003303032121)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_CQ),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_BQ),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_A5Q),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_BO5),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fb0bf000fb0b)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffef0f40f0e0004)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_BLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafff0)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y111_SLICE_X14Y111_AO6),
.Q(CLBLM_R_X11Y111_SLICE_X14Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffeeee)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_D5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_BQ),
.I5(CLBLM_R_X11Y115_SLICE_X14Y115_DQ),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffeeee)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_CLUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_CQ),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_BLUT (
.I0(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_DQ),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_D5Q),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0ac00330033)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_A5Q),
.I1(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X16Y112_DO6),
.Q(CLBLM_R_X11Y111_SLICE_X15Y111_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.Q(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y111_SLICE_X15Y111_BO6),
.Q(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_B5Q),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_DQ),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_DQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_DO6),
.I2(CLBLM_L_X12Y111_SLICE_X16Y111_CO6),
.I3(CLBLM_R_X11Y111_SLICE_X14Y111_DO6),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_CQ),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffc8ff00ffc8)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_BLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefececefefccecc)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_ALUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_C5Q),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X14Y112_AO6),
.Q(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X14Y112_BO6),
.Q(CLBLM_R_X11Y112_SLICE_X14Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X14Y112_CO6),
.Q(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X14Y112_DO6),
.Q(CLBLM_R_X11Y112_SLICE_X14Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000faff0a0f)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_DLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_DO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff411400004114)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_AQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y112_SLICE_X16Y112_A5Q),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_CO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055440000)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_BQ),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_CQ),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_BO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00bebeff00bebe)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_ALUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I1(CLBLM_R_X11Y112_SLICE_X15Y112_DO6),
.I2(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_AO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X15Y112_AO6),
.Q(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.Q(CLBLM_R_X11Y112_SLICE_X15Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000003000000010)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_DLUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I1(CLBLM_L_X12Y112_SLICE_X16Y112_BQ),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I3(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.I4(CLBLM_L_X12Y112_SLICE_X17Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c5c5c0c0c0c0)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_CO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cac000ff55ff)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_BLUT (
.I0(CLBLM_L_X12Y113_SLICE_X17Y113_CQ),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_BO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afa003030000)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_ALUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_CQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_AO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_BO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_CO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbffffffff)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_AQ),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CQ),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0e4a0e4a0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_DQ),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0cfcfc0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54fe54aa00)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_CO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_AO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_BO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_DO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff00a8a8)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_DQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e0e0e0e0e0e0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_CLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05544f0f05544)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3333aaaa3030)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_ALUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_DQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.R(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f000e0e0e0e)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_DLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_BQ),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_DQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaca0a0ffcc0000)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_CLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf088aaaa8888)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_D5Q),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30ec20f0f0a0a0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_ALUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_C5Q),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X15Y114_AO6),
.Q(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X15Y114_BO6),
.Q(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X15Y114_CO6),
.Q(CLBLM_R_X11Y114_SLICE_X15Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X15Y114_DO6),
.Q(CLBLM_R_X11Y114_SLICE_X15Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888bbb88888)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_DQ),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdce0102cdce0102)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I4(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff4400440044)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_BLUT (
.I0(CLBLM_L_X12Y115_SLICE_X16Y115_AO6),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_DQ),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0eeeeeeee)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_ALUT (
.I0(CLBLM_L_X12Y115_SLICE_X16Y115_AO6),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_BO5),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_AO6),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_BO6),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_CO6),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_DO6),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f055f000f000)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_D5Q),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddccddcc11001100)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_CLUT (
.I0(CLBLM_L_X12Y115_SLICE_X16Y115_AO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003030aaaaff00)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_BLUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_AO6),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_CQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf5f00000)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_CQ),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_BO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he0f0e0f0ffffe0f0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_DLUT (
.I0(CLBLM_L_X12Y115_SLICE_X16Y115_AO6),
.I1(CLBLM_R_X13Y115_SLICE_X19Y115_BO6),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_CQ),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_CQ),
.I4(CLBLM_R_X13Y115_SLICE_X19Y115_CO6),
.I5(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f000f0e0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_CLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000044f044f0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_DQ),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb888bb8b8)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_ALUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_CO5),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.I5(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_CO5),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_BO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_CO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_DO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddcccc11110000)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I5(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc1100fc30fc30)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_B5Q),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_CQ),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'habab0101aeae0404)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_DQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd88888fff00000)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_DQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X15Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X15Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X15Y116_BO6),
.Q(CLBLM_R_X11Y116_SLICE_X15Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X15Y116_CO6),
.Q(CLBLM_R_X11Y116_SLICE_X15Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00bfffff33000000)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_DLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_CO5),
.I1(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5b1b1e4e4a0a0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_DO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaffaaee)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I1(CLBLM_R_X11Y116_SLICE_X15Y116_BQ),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff030003ff210021)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_ALUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_DO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I5(CLBLM_L_X12Y117_SLICE_X16Y117_CO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_BO5),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_BO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00c00000ff3f)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_DO6),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h08a8882808a8882a)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_CLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafaaaffffcc00)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_CO6),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44ff040f44ff040f)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_AO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_BO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f5f0f5f0f0f0f0f)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_DLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CQ),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000232300003330)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_CLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_BO5),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeff0455aeaa0400)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.I2(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I5(CLBLM_L_X12Y114_SLICE_X17Y114_CQ),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff541000005410)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_CO6),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_B5Q),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_CO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_BO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808088810101000)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_DLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I5(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff000000cfcf)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c0f0f000ccffff)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I2(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_DO6),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8400cccca500ffff)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcddc3223cccc3333)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.I4(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3323323333333333)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.I4(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8acf0a0f2a3f0a0f)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_BLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I5(CLBLM_R_X11Y118_SLICE_X15Y118_CO6),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0f00005f0f5f0f)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_ALUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_DO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.Q(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00b8003000300030)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_DLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.I5(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc39cc39cc39cc33)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_CLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_BO6),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088880000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I1(CLBLM_L_X12Y118_SLICE_X16Y118_AO6),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303333f030ff33)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_A5Q),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_CO6),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_AO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00f0fa587)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_BLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I1(CLBLM_L_X12Y118_SLICE_X16Y118_AO5),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I3(CLBLM_L_X12Y118_SLICE_X16Y118_AO6),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcf00000fcf0fcf)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacfc0cfc0c)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I1(RIOB33_X105Y125_IOB_X1Y126_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X17Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y108_SLICE_X18Y108_AO6),
.Q(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_DO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_CO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_BO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000cf0ff000f)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_CO6),
.I4(CLBLM_R_X13Y109_SLICE_X18Y109_DQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_AO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_DO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_CO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_BO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_AO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y109_SLICE_X18Y109_AO6),
.Q(CLBLM_R_X13Y109_SLICE_X18Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y109_SLICE_X18Y109_BO6),
.Q(CLBLM_R_X13Y109_SLICE_X18Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y109_SLICE_X18Y109_CO6),
.Q(CLBLM_R_X13Y109_SLICE_X18Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y109_SLICE_X18Y109_DO6),
.Q(CLBLM_R_X13Y109_SLICE_X18Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccccf0a0)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_D5Q),
.I2(CLBLM_R_X13Y109_SLICE_X18Y109_DQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_DO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffccffaaffc0)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_CLUT (
.I0(CLBLM_R_X13Y115_SLICE_X19Y115_AQ),
.I1(CLBLM_R_X13Y109_SLICE_X18Y109_CQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_CO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4a0f5a0a0a0f5)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y109_SLICE_X18Y109_BQ),
.I2(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I3(CLBLM_L_X12Y109_SLICE_X17Y109_CO6),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_BO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf333aaaac000)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_ALUT (
.I0(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I2(CLBLM_R_X13Y109_SLICE_X18Y109_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_AO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_DO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_CO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_BO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_AO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y110_SLICE_X18Y110_AO6),
.Q(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_DO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_CO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_BO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff3f00000f3f0)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I2(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_A5Q),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_AO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_DO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_CO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_BO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_AO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y111_SLICE_X18Y111_AO6),
.Q(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y111_SLICE_X18Y111_BO6),
.Q(CLBLM_R_X13Y111_SLICE_X18Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y111_SLICE_X18Y111_CO6),
.Q(CLBLM_R_X13Y111_SLICE_X18Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h020a0000070f0000)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_DLUT (
.I0(CLBLM_R_X13Y111_SLICE_X19Y111_AQ),
.I1(CLBLM_R_X13Y111_SLICE_X19Y111_BQ),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_BQ),
.I4(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_DO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaa0500aeaa0400)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I5(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_CO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeaaaaeccca000)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_BLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_AO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y111_SLICE_X18Y111_DO6),
.I3(CLBLM_R_X13Y111_SLICE_X19Y111_BQ),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_CQ),
.I5(CLBLM_R_X13Y111_SLICE_X18Y111_BQ),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8ffa2a8a8a2a2)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_ALUT (
.I0(CLBLM_L_X12Y118_SLICE_X16Y118_BO6),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I2(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y111_SLICE_X17Y111_DO6),
.I5(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_AO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.Q(CLBLM_R_X13Y111_SLICE_X19Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y111_SLICE_X19Y111_BO6),
.Q(CLBLM_R_X13Y111_SLICE_X19Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_DO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_CO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f0f4f001000400)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I1(CLBLM_R_X13Y111_SLICE_X19Y111_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_DO6),
.I5(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_BO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff140014ff000000)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_ALUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_DO5),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_AO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y112_SLICE_X18Y112_AO6),
.Q(CLBLM_R_X13Y112_SLICE_X18Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_DO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_CO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_BO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff0000330000)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_AO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y112_SLICE_X19Y112_AO5),
.Q(CLBLM_R_X13Y112_SLICE_X19Y112_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y112_SLICE_X19Y112_BO5),
.Q(CLBLM_R_X13Y112_SLICE_X19Y112_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.Q(CLBLM_R_X13Y112_SLICE_X19Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y112_SLICE_X19Y112_BO6),
.Q(CLBLM_R_X13Y112_SLICE_X19Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_DO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_CO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc33aa99aaaa)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_BLUT (
.I0(CLBLM_R_X13Y112_SLICE_X19Y112_B5Q),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y115_SLICE_X16Y115_CO6),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_BO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111000000ffff00)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_ALUT (
.I0(CLBLM_R_X13Y112_SLICE_X19Y112_B5Q),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y115_SLICE_X16Y115_CO6),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_AO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y113_SLICE_X18Y113_AO6),
.Q(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_DO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_CO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_BO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fffc00f000fc)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_AO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_DO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_CO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_AO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y114_SLICE_X18Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y114_SLICE_X18Y114_AO6),
.Q(CLBLM_R_X13Y114_SLICE_X18Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y114_SLICE_X18Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X18Y114_DO5),
.O6(CLBLM_R_X13Y114_SLICE_X18Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y114_SLICE_X18Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X18Y114_CO5),
.O6(CLBLM_R_X13Y114_SLICE_X18Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y114_SLICE_X18Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X18Y114_BO5),
.O6(CLBLM_R_X13Y114_SLICE_X18Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00f0aaaa)
  ) CLBLM_R_X13Y114_SLICE_X18Y114_ALUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_DQ),
.I2(CLBLM_R_X13Y114_SLICE_X18Y114_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y114_SLICE_X18Y114_AO5),
.O6(CLBLM_R_X13Y114_SLICE_X18Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y114_SLICE_X19Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X19Y114_DO5),
.O6(CLBLM_R_X13Y114_SLICE_X19Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y114_SLICE_X19Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X19Y114_CO5),
.O6(CLBLM_R_X13Y114_SLICE_X19Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y114_SLICE_X19Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X19Y114_BO5),
.O6(CLBLM_R_X13Y114_SLICE_X19Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y114_SLICE_X19Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X19Y114_AO5),
.O6(CLBLM_R_X13Y114_SLICE_X19Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y115_SLICE_X18Y115_AO6),
.Q(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y115_SLICE_X18Y115_BO6),
.Q(CLBLM_R_X13Y115_SLICE_X18Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_DO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808101008881000)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_CLUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I1(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I4(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I5(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_CO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fcf0fd000c000d)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I1(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_BO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00fc00cf)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_ALUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I1(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.I2(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I3(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_AO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X13Y114_SLICE_X18Y114_AQ),
.Q(CLBLM_R_X13Y115_SLICE_X19Y115_AQ),
.R(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00000000)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_DLUT (
.I0(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y116_SLICE_X15Y116_A5Q),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_DO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0000000f00)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_CO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7531dfdf2f2fd0d0)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I4(CLBLM_R_X13Y115_SLICE_X19Y115_DO6),
.I5(CLBLM_R_X13Y115_SLICE_X19Y115_AO5),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_BO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2020202005050f0f)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_AO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y116_SLICE_X18Y116_AO6),
.Q(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y116_SLICE_X18Y116_BO6),
.Q(CLBLM_R_X13Y116_SLICE_X18Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X18Y116_DO5),
.O6(CLBLM_R_X13Y116_SLICE_X18Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X18Y116_CO5),
.O6(CLBLM_R_X13Y116_SLICE_X18Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4f5f5a0e4a0a0)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y116_SLICE_X18Y116_BQ),
.I2(CLBLM_R_X13Y112_SLICE_X18Y112_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.I5(CLBLM_R_X11Y116_SLICE_X15Y116_BQ),
.O5(CLBLM_R_X13Y116_SLICE_X18Y116_BO5),
.O6(CLBLM_R_X13Y116_SLICE_X18Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaac0f0)
  ) CLBLM_R_X13Y116_SLICE_X18Y116_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.I2(CLBLM_R_X13Y116_SLICE_X18Y116_AQ),
.I3(CLBLM_R_X13Y117_SLICE_X18Y117_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y117_SLICE_X16Y117_CO6),
.O5(CLBLM_R_X13Y116_SLICE_X18Y116_AO5),
.O6(CLBLM_R_X13Y116_SLICE_X18Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X19Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X19Y116_DO5),
.O6(CLBLM_R_X13Y116_SLICE_X19Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X19Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X19Y116_CO5),
.O6(CLBLM_R_X13Y116_SLICE_X19Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X19Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X19Y116_BO5),
.O6(CLBLM_R_X13Y116_SLICE_X19Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y116_SLICE_X19Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y116_SLICE_X19Y116_AO5),
.O6(CLBLM_R_X13Y116_SLICE_X19Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y117_SLICE_X18Y117_AO6),
.Q(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100010001000000)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_DLUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I1(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I5(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_DO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_CLUT (
.I0(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.I1(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.I2(CLBLM_L_X12Y113_SLICE_X17Y113_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I4(CLBLM_R_X13Y117_SLICE_X18Y117_DO6),
.I5(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_CO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50500003af23cc30)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f2f203030202)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_ALUT (
.I0(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y118_SLICE_X17Y118_AO6),
.I5(CLBLM_L_X12Y112_SLICE_X17Y112_CQ),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_AO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_DO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_CO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_BO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_AO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y118_SLICE_X18Y118_AO6),
.Q(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_DO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_CO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_BO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0fcf0fc)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I4(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_AO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_DO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_CO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_BO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_AO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y115_SLICE_X56Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y115_SLICE_X56Y115_DO5),
.O6(CLBLM_R_X37Y115_SLICE_X56Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y115_SLICE_X56Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y115_SLICE_X56Y115_CO5),
.O6(CLBLM_R_X37Y115_SLICE_X56Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y115_SLICE_X56Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y115_SLICE_X56Y115_BO5),
.O6(CLBLM_R_X37Y115_SLICE_X56Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000505000005050)
  ) CLBLM_R_X37Y115_SLICE_X56Y115_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(1'b1),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.I5(1'b1),
.O5(CLBLM_R_X37Y115_SLICE_X56Y115_AO5),
.O6(CLBLM_R_X37Y115_SLICE_X56Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y115_SLICE_X57Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y115_SLICE_X57Y115_DO5),
.O6(CLBLM_R_X37Y115_SLICE_X57Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y115_SLICE_X57Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y115_SLICE_X57Y115_CO5),
.O6(CLBLM_R_X37Y115_SLICE_X57Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y115_SLICE_X57Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y115_SLICE_X57Y115_BO5),
.O6(CLBLM_R_X37Y115_SLICE_X57Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y115_SLICE_X57Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y115_SLICE_X57Y115_AO5),
.O6(CLBLM_R_X37Y115_SLICE_X57Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_ALUT (
.I0(RIOB33_X105Y139_IOB_X1Y139_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfffff0f0ffff)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555f5f5f5f5)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffaaaaffff)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_ALUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafafffffafa)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(1'b1),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(1'b1),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555f5f5f5f5)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(1'b1),
.I2(CLBLM_R_X13Y115_SLICE_X19Y115_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_CO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_AO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_DO6),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_L_X12Y110_SLICE_X16Y110_D5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_L_X12Y110_SLICE_X16Y110_DQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X4Y112_SLICE_X5Y112_CQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X10Y111_SLICE_X12Y111_DQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_R_X11Y120_SLICE_X14Y120_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X7Y117_SLICE_X8Y117_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_L_X8Y113_SLICE_X10Y113_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X4Y112_SLICE_X5Y112_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_L_X10Y115_SLICE_X12Y115_D5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X4Y112_SLICE_X5Y112_BQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_L_X8Y123_SLICE_X11Y123_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X7Y119_SLICE_X8Y119_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y138_SLICE_X163Y138_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_L_X8Y150_SLICE_X10Y150_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_BO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLM_R_X37Y115_SLICE_X56Y115_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_L_X12Y112_SLICE_X17Y112_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_L_X12Y112_SLICE_X17Y112_DO5),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X8Y150_SLICE_X10Y150_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO6),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_L_X10Y122_SLICE_X12Y122_BO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_L_X12Y122_SLICE_X17Y122_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_L_X12Y112_SLICE_X17Y112_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_L_X12Y112_SLICE_X17Y112_DO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X13Y118_SLICE_X18Y118_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_R_X13Y115_SLICE_X19Y115_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y118_SLICE_X17Y118_AQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_BO6),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_BO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_AMUX = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_BMUX = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_CMUX = CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_DMUX = CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_AMUX = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_AMUX = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_CMUX = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_AMUX = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_AMUX = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_AMUX = CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_BMUX = CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_CMUX = CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_AMUX = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_BMUX = CLBLL_L_X4Y108_SLICE_X4Y108_B5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_CMUX = CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_AMUX = CLBLL_L_X4Y109_SLICE_X5Y109_A5Q;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_CMUX = CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_CMUX = CLBLL_L_X4Y110_SLICE_X4Y110_C5Q;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_BMUX = CLBLL_L_X4Y110_SLICE_X5Y110_B5Q;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_DMUX = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_CMUX = CLBLL_L_X4Y112_SLICE_X5Y112_C5Q;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_CMUX = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_CMUX = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_AMUX = CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_BMUX = CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CMUX = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_AMUX = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_DMUX = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_AMUX = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_BMUX = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_DMUX = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_AMUX = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_AMUX = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_BMUX = CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_AMUX = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_AMUX = CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_BMUX = CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_DMUX = CLBLM_L_X8Y107_SLICE_X10Y107_DO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_AMUX = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_DMUX = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_DMUX = CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_AMUX = CLBLM_L_X8Y109_SLICE_X11Y109_A5Q;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_DMUX = CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_DMUX = CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_CMUX = CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_AMUX = CLBLM_L_X8Y111_SLICE_X10Y111_A5Q;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_BMUX = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_CMUX = CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_CMUX = CLBLM_L_X8Y113_SLICE_X10Y113_C5Q;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_CMUX = CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_DMUX = CLBLM_L_X8Y114_SLICE_X10Y114_D5Q;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_AMUX = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_DMUX = CLBLM_L_X8Y115_SLICE_X10Y115_DO5;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_BMUX = CLBLM_L_X8Y115_SLICE_X11Y115_B5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_AMUX = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_CMUX = CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A = CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B = CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B = CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_AMUX = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_AMUX = CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_CMUX = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A = CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B = CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C = CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A = CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A = CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_AMUX = CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A = CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C = CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_CMUX = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_AMUX = CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_DMUX = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_AMUX = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_CMUX = CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_DMUX = CLBLM_L_X10Y111_SLICE_X12Y111_D5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_BMUX = CLBLM_L_X10Y111_SLICE_X13Y111_B5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_CMUX = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_DMUX = CLBLM_L_X10Y111_SLICE_X13Y111_D5Q;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_BMUX = CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_DMUX = CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_DMUX = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_AMUX = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_AMUX = CLBLM_L_X10Y114_SLICE_X13Y114_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_CMUX = CLBLM_L_X10Y114_SLICE_X13Y114_C5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B = CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C = CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D = CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_CMUX = CLBLM_L_X10Y115_SLICE_X12Y115_C5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_DMUX = CLBLM_L_X10Y115_SLICE_X12Y115_D5Q;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A = CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B = CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_CMUX = CLBLM_L_X10Y116_SLICE_X12Y116_C5Q;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_DMUX = CLBLM_L_X10Y116_SLICE_X12Y116_D5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A = CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_AMUX = CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A = CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_BMUX = CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_CMUX = CLBLM_L_X10Y118_SLICE_X12Y118_C5Q;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_AMUX = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_BMUX = CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_AMUX = CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_BMUX = CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_CMUX = CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_AMUX = CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_BMUX = CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A = CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_AMUX = CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_DMUX = CLBLM_L_X12Y107_SLICE_X16Y107_DO5;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C = CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_BMUX = CLBLM_L_X12Y109_SLICE_X16Y109_BO5;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_CMUX = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_DMUX = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D = CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_DMUX = CLBLM_L_X12Y110_SLICE_X16Y110_D5Q;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A = CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B = CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C = CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D = CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_BMUX = CLBLM_L_X12Y111_SLICE_X16Y111_B5Q;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A = CLBLM_L_X12Y111_SLICE_X17Y111_AO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B = CLBLM_L_X12Y111_SLICE_X17Y111_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C = CLBLM_L_X12Y111_SLICE_X17Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D = CLBLM_L_X12Y111_SLICE_X17Y111_DO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_CMUX = CLBLM_L_X12Y111_SLICE_X17Y111_CO5;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A = CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B = CLBLM_L_X12Y112_SLICE_X16Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C = CLBLM_L_X12Y112_SLICE_X16Y112_CO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D = CLBLM_L_X12Y112_SLICE_X16Y112_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_AMUX = CLBLM_L_X12Y112_SLICE_X16Y112_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_BMUX = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_CMUX = CLBLM_L_X12Y112_SLICE_X16Y112_CO5;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_DMUX = CLBLM_L_X12Y112_SLICE_X16Y112_DO5;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A = CLBLM_L_X12Y112_SLICE_X17Y112_AO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B = CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C = CLBLM_L_X12Y112_SLICE_X17Y112_CO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_DMUX = CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A = CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C = CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D = CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A = CLBLM_L_X12Y113_SLICE_X17Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B = CLBLM_L_X12Y113_SLICE_X17Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C = CLBLM_L_X12Y113_SLICE_X17Y113_CO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D = CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A = CLBLM_L_X12Y114_SLICE_X16Y114_AO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A = CLBLM_L_X12Y114_SLICE_X17Y114_AO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B = CLBLM_L_X12Y114_SLICE_X17Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C = CLBLM_L_X12Y114_SLICE_X17Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D = CLBLM_L_X12Y114_SLICE_X17Y114_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_AMUX = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_DMUX = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A = CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B = CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C = CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_DMUX = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A = CLBLM_L_X12Y116_SLICE_X16Y116_AO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B = CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D = CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_BMUX = CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_CMUX = CLBLM_L_X12Y116_SLICE_X16Y116_CO5;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A = CLBLM_L_X12Y116_SLICE_X17Y116_AO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B = CLBLM_L_X12Y116_SLICE_X17Y116_BO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C = CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D = CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_CMUX = CLBLM_L_X12Y116_SLICE_X17Y116_CO5;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C = CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D = CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_BMUX = CLBLM_L_X12Y117_SLICE_X16Y117_BO5;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_CMUX = CLBLM_L_X12Y117_SLICE_X16Y117_CO5;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A = CLBLM_L_X12Y117_SLICE_X17Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B = CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D = CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A = CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C = CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D = CLBLM_L_X12Y118_SLICE_X16Y118_DO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_AMUX = CLBLM_L_X12Y118_SLICE_X16Y118_AO5;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A = CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B = CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C = CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A = CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B = CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A = CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_AMUX = CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_CMUX = CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_DMUX = CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_CMUX = CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_CMUX = CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_DMUX = CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_DMUX = CLBLM_R_X3Y110_SLICE_X3Y110_D5Q;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_AMUX = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_AMUX = CLBLM_R_X3Y111_SLICE_X3Y111_A5Q;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_DMUX = CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_BMUX = CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_CMUX = CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_DMUX = CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_AMUX = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_AMUX = CLBLM_R_X3Y114_SLICE_X2Y114_A5Q;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_AMUX = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_DMUX = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_DMUX = CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_BMUX = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_CMUX = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_DMUX = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_CMUX = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_AMUX = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_AMUX = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_BMUX = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_DMUX = CLBLM_R_X5Y107_SLICE_X7Y107_D5Q;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_AMUX = CLBLM_R_X5Y109_SLICE_X7Y109_A5Q;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_BMUX = CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_CMUX = CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_DMUX = CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_CMUX = CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_AMUX = CLBLM_R_X5Y112_SLICE_X7Y112_A5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_BMUX = CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_DMUX = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_BMUX = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_AMUX = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_DMUX = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_AMUX = CLBLM_R_X5Y116_SLICE_X6Y116_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CMUX = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_DMUX = CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_BMUX = CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_CMUX = CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_AMUX = CLBLM_R_X5Y117_SLICE_X7Y117_A5Q;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_AMUX = CLBLM_R_X5Y119_SLICE_X6Y119_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_BMUX = CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CMUX = CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A = CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B = CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A = CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B = CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_BMUX = CLBLM_R_X7Y106_SLICE_X9Y106_B5Q;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_CMUX = CLBLM_R_X7Y107_SLICE_X8Y107_CO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_AMUX = CLBLM_R_X7Y107_SLICE_X9Y107_A5Q;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_BMUX = CLBLM_R_X7Y107_SLICE_X9Y107_B5Q;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_CMUX = CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_BMUX = CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_DMUX = CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_AMUX = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_CMUX = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_DMUX = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_CMUX = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_BMUX = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_DMUX = CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_AMUX = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_AMUX = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_BMUX = CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_BMUX = CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_CMUX = CLBLM_R_X7Y114_SLICE_X8Y114_C5Q;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_DMUX = CLBLM_R_X7Y114_SLICE_X8Y114_D5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_CMUX = CLBLM_R_X7Y114_SLICE_X9Y114_C5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_DMUX = CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_AMUX = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_CMUX = CLBLM_R_X7Y116_SLICE_X8Y116_C5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_BMUX = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_AMUX = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_DMUX = CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_AMUX = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_CMUX = CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B = CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_BMUX = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_AMUX = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_BMUX = CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_DMUX = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_AMUX = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_BMUX = CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_CMUX = CLBLM_R_X11Y107_SLICE_X14Y107_CO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_CMUX = CLBLM_R_X11Y107_SLICE_X15Y107_CO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_DMUX = CLBLM_R_X11Y107_SLICE_X15Y107_DO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_BMUX = CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_AMUX = CLBLM_R_X11Y109_SLICE_X14Y109_A5Q;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_BMUX = CLBLM_R_X11Y109_SLICE_X14Y109_BO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_AMUX = CLBLM_R_X11Y110_SLICE_X14Y110_A5Q;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_AMUX = CLBLM_R_X11Y110_SLICE_X15Y110_A5Q;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_AMUX = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_AMUX = CLBLM_R_X11Y111_SLICE_X15Y111_A5Q;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_CMUX = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_DMUX = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C = CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D = CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A = CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_AMUX = CLBLM_R_X11Y112_SLICE_X15Y112_AO5;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_BMUX = CLBLM_R_X11Y112_SLICE_X15Y112_BO5;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_DMUX = CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B = CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_AMUX = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_CMUX = CLBLM_R_X11Y113_SLICE_X15Y113_CO5;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_AMUX = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_BMUX = CLBLM_R_X11Y114_SLICE_X14Y114_BO5;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_CMUX = CLBLM_R_X11Y114_SLICE_X14Y114_CO5;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_DMUX = CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D = CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_BMUX = CLBLM_R_X11Y115_SLICE_X14Y115_B5Q;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A = CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_AMUX = CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_CMUX = CLBLM_R_X11Y116_SLICE_X14Y116_C5Q;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_AMUX = CLBLM_R_X11Y116_SLICE_X15Y116_A5Q;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_DMUX = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_BMUX = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_CMUX = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A = CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A = CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B = CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C = CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_AMUX = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_CMUX = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_DMUX = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A = CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_BMUX = CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_AMUX = CLBLM_R_X11Y120_SLICE_X14Y120_A5Q;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A = CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B = CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C = CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A = CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A = CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D = CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A = CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B = CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C = CLBLM_R_X13Y108_SLICE_X19Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D = CLBLM_R_X13Y108_SLICE_X19Y108_DO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A = CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B = CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C = CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D = CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A = CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B = CLBLM_R_X13Y109_SLICE_X19Y109_BO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C = CLBLM_R_X13Y109_SLICE_X19Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D = CLBLM_R_X13Y109_SLICE_X19Y109_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A = CLBLM_R_X13Y110_SLICE_X18Y110_AO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B = CLBLM_R_X13Y110_SLICE_X18Y110_BO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C = CLBLM_R_X13Y110_SLICE_X18Y110_CO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A = CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B = CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C = CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D = CLBLM_R_X13Y110_SLICE_X19Y110_DO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A = CLBLM_R_X13Y111_SLICE_X18Y111_AO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B = CLBLM_R_X13Y111_SLICE_X18Y111_BO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C = CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_DMUX = CLBLM_R_X13Y111_SLICE_X18Y111_DO5;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B = CLBLM_R_X13Y111_SLICE_X19Y111_BO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C = CLBLM_R_X13Y111_SLICE_X19Y111_CO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D = CLBLM_R_X13Y111_SLICE_X19Y111_DO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A = CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B = CLBLM_R_X13Y112_SLICE_X18Y112_BO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C = CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D = CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B = CLBLM_R_X13Y112_SLICE_X19Y112_BO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C = CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_AMUX = CLBLM_R_X13Y112_SLICE_X19Y112_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_BMUX = CLBLM_R_X13Y112_SLICE_X19Y112_B5Q;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A = CLBLM_R_X13Y113_SLICE_X18Y113_AO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B = CLBLM_R_X13Y113_SLICE_X18Y113_BO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C = CLBLM_R_X13Y113_SLICE_X18Y113_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D = CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A = CLBLM_R_X13Y113_SLICE_X19Y113_AO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B = CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D = CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A = CLBLM_R_X13Y114_SLICE_X18Y114_AO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B = CLBLM_R_X13Y114_SLICE_X18Y114_BO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C = CLBLM_R_X13Y114_SLICE_X18Y114_CO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D = CLBLM_R_X13Y114_SLICE_X18Y114_DO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A = CLBLM_R_X13Y114_SLICE_X19Y114_AO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C = CLBLM_R_X13Y114_SLICE_X19Y114_CO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D = CLBLM_R_X13Y114_SLICE_X19Y114_DO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A = CLBLM_R_X13Y115_SLICE_X18Y115_AO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B = CLBLM_R_X13Y115_SLICE_X18Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C = CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D = CLBLM_R_X13Y115_SLICE_X18Y115_DO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A = CLBLM_R_X13Y115_SLICE_X19Y115_AO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B = CLBLM_R_X13Y115_SLICE_X19Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C = CLBLM_R_X13Y115_SLICE_X19Y115_CO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D = CLBLM_R_X13Y115_SLICE_X19Y115_DO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_AMUX = CLBLM_R_X13Y115_SLICE_X19Y115_AO5;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A = CLBLM_R_X13Y116_SLICE_X18Y116_AO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B = CLBLM_R_X13Y116_SLICE_X18Y116_BO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C = CLBLM_R_X13Y116_SLICE_X18Y116_CO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D = CLBLM_R_X13Y116_SLICE_X18Y116_DO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A = CLBLM_R_X13Y116_SLICE_X19Y116_AO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B = CLBLM_R_X13Y116_SLICE_X19Y116_BO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C = CLBLM_R_X13Y116_SLICE_X19Y116_CO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D = CLBLM_R_X13Y116_SLICE_X19Y116_DO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A = CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B = CLBLM_R_X13Y117_SLICE_X18Y117_BO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C = CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D = CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_BMUX = CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A = CLBLM_R_X13Y117_SLICE_X19Y117_AO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B = CLBLM_R_X13Y117_SLICE_X19Y117_BO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C = CLBLM_R_X13Y117_SLICE_X19Y117_CO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D = CLBLM_R_X13Y117_SLICE_X19Y117_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A = CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B = CLBLM_R_X13Y118_SLICE_X18Y118_BO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C = CLBLM_R_X13Y118_SLICE_X18Y118_CO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D = CLBLM_R_X13Y118_SLICE_X18Y118_DO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A = CLBLM_R_X13Y118_SLICE_X19Y118_AO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B = CLBLM_R_X13Y118_SLICE_X19Y118_BO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C = CLBLM_R_X13Y118_SLICE_X19Y118_CO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D = CLBLM_R_X13Y118_SLICE_X19Y118_DO6;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_A = CLBLM_R_X37Y115_SLICE_X56Y115_AO6;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_B = CLBLM_R_X37Y115_SLICE_X56Y115_BO6;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_C = CLBLM_R_X37Y115_SLICE_X56Y115_CO6;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_D = CLBLM_R_X37Y115_SLICE_X56Y115_DO6;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_A = CLBLM_R_X37Y115_SLICE_X57Y115_AO6;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_B = CLBLM_R_X37Y115_SLICE_X57Y115_BO6;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_C = CLBLM_R_X37Y115_SLICE_X57Y115_CO6;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_D = CLBLM_R_X37Y115_SLICE_X57Y115_DO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A = CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B = CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C = CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D = CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B = CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C = CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D = CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_AMUX = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A = CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B = CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C = CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D = CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B = CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C = CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D = CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_AMUX = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A = CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B = CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C = CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D = CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B = CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C = CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D = CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_AMUX = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_L_X12Y110_SLICE_X16Y110_D5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_L_X12Y110_SLICE_X16Y110_DQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X4Y112_SLICE_X5Y112_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_R_X11Y120_SLICE_X14Y120_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X4Y112_SLICE_X5Y112_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_L_X8Y113_SLICE_X10Y113_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_L_X10Y115_SLICE_X12Y115_D5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X4Y112_SLICE_X5Y112_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X10Y111_SLICE_X12Y111_DQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y118_SLICE_X17Y118_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_R_X13Y115_SLICE_X19Y115_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLM_R_X37Y115_SLICE_X56Y115_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = CLBLM_R_X7Y108_SLICE_X8Y108_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = 1'b1;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = CLBLM_R_X3Y110_SLICE_X3Y110_D5Q;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A1 = CLBLM_L_X12Y114_SLICE_X17Y114_DO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A2 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A3 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A6 = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B2 = CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B3 = CLBLM_R_X7Y106_SLICE_X8Y106_BQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B4 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B5 = CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B6 = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLM_R_X37Y115_SLICE_X56Y115_AO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C1 = CLBLM_R_X13Y114_SLICE_X18Y114_AQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C2 = CLBLM_L_X12Y114_SLICE_X17Y114_CQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C3 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C5 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C6 = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D1 = CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D2 = CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D3 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D4 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D5 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D6 = CLBLM_L_X12Y114_SLICE_X16Y114_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A1 = CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A4 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A6 = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B1 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B2 = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B3 = CLBLM_L_X12Y114_SLICE_X16Y114_CQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B5 = CLBLM_L_X12Y114_SLICE_X16Y114_BQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C2 = CLBLM_L_X12Y114_SLICE_X16Y114_CQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C3 = CLBLM_R_X13Y116_SLICE_X18Y116_BQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C4 = CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C5 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C6 = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = 1'b1;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_BQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D3 = CLBLM_L_X12Y114_SLICE_X16Y114_DQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D4 = CLBLM_R_X11Y114_SLICE_X15Y114_DQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D5 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D6 = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A2 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B2 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C2 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D2 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A2 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A4 = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A5 = CLBLM_R_X13Y109_SLICE_X18Y109_DQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B2 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C2 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D2 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A1 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A1 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A2 = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A3 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A4 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A5 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A6 = CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B1 = CLBLM_R_X13Y114_SLICE_X18Y114_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B2 = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B3 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B4 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B5 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B6 = CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C1 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C2 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C3 = CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C4 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C5 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D1 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D2 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D3 = CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D4 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D5 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D6 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A1 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A2 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A4 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A5 = CLBLM_L_X12Y116_SLICE_X17Y116_CO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_AX = CLBLM_L_X12Y110_SLICE_X16Y110_DQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B1 = CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B2 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B3 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B4 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B5 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B6 = CLBLM_L_X12Y114_SLICE_X16Y114_CQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A2 = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C1 = CLBLM_L_X12Y116_SLICE_X17Y116_CO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C2 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C3 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C5 = CLBLM_R_X13Y115_SLICE_X19Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C6 = CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D2 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D3 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D4 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D5 = CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_SR = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A1 = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A2 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A3 = CLBLM_R_X13Y109_SLICE_X18Y109_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A6 = CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B2 = CLBLM_R_X13Y109_SLICE_X18Y109_BQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B3 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B4 = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B5 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C1 = CLBLM_R_X13Y115_SLICE_X19Y115_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C2 = CLBLM_R_X13Y109_SLICE_X18Y109_CQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C4 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D2 = CLBLM_L_X10Y111_SLICE_X13Y111_D5Q;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D3 = CLBLM_R_X13Y109_SLICE_X18Y109_DQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D6 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C1 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C2 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C4 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_C6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A1 = CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A2 = CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A3 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A5 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A6 = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B1 = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B2 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B5 = CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B6 = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A1 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A2 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A3 = CLBLM_R_X7Y106_SLICE_X9Y106_B5Q;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A4 = CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_DQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A6 = CLBLM_L_X10Y107_SLICE_X13Y107_CQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C1 = CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C2 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B1 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B2 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B4 = CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_DQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B6 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D1 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C1 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C4 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C6 = CLBLM_L_X10Y106_SLICE_X12Y106_BQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D3 = CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D4 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D5 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D6 = CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A1 = CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A3 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D1 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D2 = CLBLM_R_X11Y111_SLICE_X15Y111_A5Q;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D3 = CLBLM_R_X5Y107_SLICE_X7Y107_D5Q;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D4 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D6 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B1 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B3 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A1 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A5 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A6 = CLBLM_L_X10Y114_SLICE_X12Y114_CQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C1 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C2 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B3 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B4 = CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B5 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B6 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D1 = CLBLM_R_X11Y116_SLICE_X15Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D2 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C1 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C2 = CLBLM_L_X10Y106_SLICE_X12Y106_CQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C4 = CLBLM_L_X10Y107_SLICE_X13Y107_CQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C5 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D3 = CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D4 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D6 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A3 = CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A4 = CLBLM_R_X13Y117_SLICE_X18Y117_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D1 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D2 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D4 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_A6 = CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C4 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C5 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B2 = CLBLM_R_X13Y116_SLICE_X18Y116_BQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B3 = CLBLM_R_X13Y112_SLICE_X18Y112_AQ;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B4 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B5 = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B6 = CLBLM_R_X11Y116_SLICE_X15Y116_BQ;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D6 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A2 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A3 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D1 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A6 = CLBLM_R_X11Y110_SLICE_X14Y110_A5Q;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B3 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D3 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D4 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C2 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D5 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D6 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C6 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A3 = CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A4 = CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A5 = CLBLM_L_X10Y109_SLICE_X13Y109_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A6 = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B1 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B2 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B3 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B4 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B5 = CLBLM_R_X13Y116_SLICE_X18Y116_BQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B6 = CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B3 = CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B4 = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A1 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A2 = CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A3 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A4 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A5 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C1 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C2 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B1 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B2 = CLBLM_L_X10Y107_SLICE_X13Y107_BQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B3 = CLBLM_L_X10Y109_SLICE_X13Y109_BQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B5 = CLBLM_R_X11Y116_SLICE_X14Y116_DQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D2 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C1 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C2 = CLBLM_L_X10Y107_SLICE_X13Y107_CQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C3 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C4 = CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C5 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D3 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D4 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D6 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A3 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A5 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D1 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D2 = CLBLM_R_X11Y110_SLICE_X14Y110_A5Q;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D3 = CLBLM_L_X10Y111_SLICE_X13Y111_CQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D4 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D5 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D6 = CLBLM_R_X11Y107_SLICE_X14Y107_CO5;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B2 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B5 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B1 = CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A3 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A4 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A5 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A6 = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C1 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C2 = CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C3 = CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B1 = CLBLM_L_X10Y109_SLICE_X13Y109_BQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B2 = CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B3 = CLBLM_L_X10Y107_SLICE_X12Y107_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B4 = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B5 = CLBLM_R_X5Y107_SLICE_X7Y107_D5Q;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D1 = CLBLM_L_X12Y117_SLICE_X16Y117_CO5;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D2 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C1 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C2 = CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C3 = CLBLM_L_X10Y111_SLICE_X13Y111_CQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C4 = CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C5 = CLBLM_L_X8Y107_SLICE_X11Y107_DQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C6 = CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D3 = CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D4 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D5 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D6 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D1 = CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D2 = CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D4 = CLBLM_L_X10Y107_SLICE_X13Y107_CQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D5 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D6 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A1 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A2 = CLBLM_R_X13Y111_SLICE_X18Y111_DO5;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A3 = CLBLM_R_X13Y111_SLICE_X19Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A5 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B2 = CLBLM_R_X13Y111_SLICE_X19Y111_BQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D5 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B5 = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B6 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C1 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C2 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C4 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C5 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C4 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C5 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C6 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D2 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D4 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D5 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D6 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A1 = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A2 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A3 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A5 = CLBLM_L_X12Y111_SLICE_X17Y111_DO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A6 = CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B1 = CLBLM_R_X11Y112_SLICE_X15Y112_AO5;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B3 = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B4 = CLBLM_R_X13Y111_SLICE_X19Y111_BQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B5 = CLBLM_R_X13Y111_SLICE_X18Y111_CQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B6 = CLBLM_R_X13Y111_SLICE_X18Y111_BQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C2 = CLBLM_R_X13Y111_SLICE_X18Y111_CQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C5 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C6 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D1 = CLBLM_R_X13Y111_SLICE_X19Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D2 = CLBLM_R_X13Y111_SLICE_X19Y111_BQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D4 = CLBLM_R_X13Y111_SLICE_X18Y111_BQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D5 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A4 = CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A6 = CLBLM_L_X10Y107_SLICE_X13Y107_CQ;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B5 = CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A1 = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A2 = CLBLM_L_X12Y114_SLICE_X17Y114_CQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A3 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A4 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A5 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A6 = CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_AX = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B1 = CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B2 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B3 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B4 = CLBLM_L_X12Y113_SLICE_X17Y113_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B5 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B6 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A1 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A3 = CLBLM_L_X10Y108_SLICE_X13Y108_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A5 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A6 = CLBLM_L_X8Y108_SLICE_X11Y108_CQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C1 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C2 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C3 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B1 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B2 = CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B3 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B4 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B5 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B6 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C1 = CLBLM_R_X11Y110_SLICE_X15Y110_BQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C2 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C4 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C5 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D2 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D3 = CLBLM_L_X10Y111_SLICE_X13Y111_CQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D4 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D5 = CLBLM_L_X8Y109_SLICE_X11Y109_A5Q;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A1 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A4 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B2 = CLBLM_L_X10Y108_SLICE_X12Y108_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B3 = CLBLM_L_X12Y108_SLICE_X16Y108_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B5 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B6 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C5 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D1 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D3 = CLBLM_L_X10Y108_SLICE_X12Y108_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D4 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D5 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D6 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A1 = CLBLM_R_X13Y112_SLICE_X19Y112_B5Q;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A2 = CLBLM_R_X13Y112_SLICE_X19Y112_BQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A4 = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A5 = CLBLM_R_X13Y112_SLICE_X19Y112_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B1 = CLBLM_R_X13Y112_SLICE_X19Y112_B5Q;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B2 = CLBLM_R_X13Y112_SLICE_X19Y112_BQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B4 = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B5 = CLBLM_R_X13Y112_SLICE_X19Y112_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C2 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D2 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A6 = CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C2 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D2 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D6 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B3 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A1 = CLBLM_R_X11Y109_SLICE_X14Y109_A5Q;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A2 = CLBLM_R_X11Y109_SLICE_X14Y109_CQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A3 = CLBLM_L_X10Y109_SLICE_X13Y109_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B1 = CLBLM_R_X13Y109_SLICE_X18Y109_CQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B2 = CLBLM_L_X10Y109_SLICE_X13Y109_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B4 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B5 = CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C1 = CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C2 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C3 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C4 = CLBLM_R_X11Y110_SLICE_X14Y110_A5Q;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C6 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D2 = CLBLM_R_X13Y109_SLICE_X18Y109_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D3 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D4 = CLBLM_L_X8Y109_SLICE_X10Y109_CQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D5 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D6 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A2 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A3 = CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A5 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B5 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B6 = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C1 = CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C2 = CLBLM_L_X10Y106_SLICE_X12Y106_CQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C3 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C4 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C5 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C6 = CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D1 = CLBLM_L_X8Y109_SLICE_X10Y109_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D2 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D4 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D6 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A1 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C6 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A3 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A5 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A6 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D6 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A1 = CLBLM_L_X10Y107_SLICE_X12Y107_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A2 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A3 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A5 = CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C3 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B1 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B2 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B3 = CLBLM_L_X10Y110_SLICE_X13Y110_CQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B4 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B6 = CLBLM_R_X11Y116_SLICE_X14Y116_DQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C2 = CLBLM_L_X10Y110_SLICE_X13Y110_CQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_CQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C6 = CLBLM_R_X13Y109_SLICE_X18Y109_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D2 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D3 = CLBLM_L_X10Y110_SLICE_X13Y110_DQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D5 = CLBLM_L_X10Y107_SLICE_X12Y107_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D6 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A3 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A4 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A5 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B2 = CLBLL_L_X4Y108_SLICE_X5Y108_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B3 = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B4 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B5 = CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C1 = CLBLM_R_X11Y110_SLICE_X15Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C3 = CLBLM_L_X10Y110_SLICE_X12Y110_DQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D2 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D3 = CLBLM_L_X10Y110_SLICE_X12Y110_DQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D4 = CLBLM_R_X3Y108_SLICE_X2Y108_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D6 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A1 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A2 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C4 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A4 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A6 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B1 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B2 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B3 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B4 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B6 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C1 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C2 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C3 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C4 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C6 = 1'b1;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D1 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D2 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D3 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D4 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D6 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A1 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A2 = CLBLM_L_X8Y113_SLICE_X11Y113_DQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A3 = CLBLM_R_X13Y114_SLICE_X18Y114_AQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A4 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A5 = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B1 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B2 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B3 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B4 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B6 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C1 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C2 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C3 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C4 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D1 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D2 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D3 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D4 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C2 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A1 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A2 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A3 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A4 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A5 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B2 = CLBLM_R_X11Y110_SLICE_X15Y110_CQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B3 = CLBLM_R_X11Y107_SLICE_X15Y107_BQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B4 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D2 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C1 = CLBLM_L_X10Y108_SLICE_X13Y108_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_A5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C5 = CLBLM_R_X11Y115_SLICE_X14Y115_DQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D3 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D4 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D1 = CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D4 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D5 = CLBLM_L_X10Y111_SLICE_X13Y111_B5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C1 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A1 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A2 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A3 = CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A4 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A6 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C2 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B1 = CLBLM_L_X8Y112_SLICE_X10Y112_DQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B2 = CLBLM_L_X10Y111_SLICE_X12Y111_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B6 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C3 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C4 = CLBLM_L_X10Y108_SLICE_X12Y108_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C5 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A1 = CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A2 = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D3 = CLBLM_R_X11Y110_SLICE_X14Y110_CQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D4 = CLBLM_L_X8Y110_SLICE_X11Y110_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B6 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A5 = CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A6 = CLBLM_L_X12Y112_SLICE_X17Y112_CQ;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B3 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C3 = 1'b1;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A1 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A2 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A3 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A5 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_AX = CLBLM_R_X13Y114_SLICE_X18Y114_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B1 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B4 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B2 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B3 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B4 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B5 = CLBLM_R_X13Y115_SLICE_X19Y115_DO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B6 = CLBLM_R_X13Y115_SLICE_X19Y115_AO5;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B2 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C4 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C5 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B4 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B5 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D1 = CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B5 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D6 = CLBLM_R_X11Y116_SLICE_X15Y116_A5Q;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_SR = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A1 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A2 = CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A3 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A4 = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A5 = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B1 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B2 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B4 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B5 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B6 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C1 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C2 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C4 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C5 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C6 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C4 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C5 = CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C6 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A2 = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A3 = CLBLM_R_X11Y116_SLICE_X15Y116_A5Q;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A4 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D2 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A6 = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A1 = CLBLM_L_X12Y118_SLICE_X17Y118_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A2 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B3 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B4 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B5 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B6 = 1'b1;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B2 = CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A2 = CLBLM_L_X10Y112_SLICE_X13Y112_DQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A3 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A6 = CLBLM_R_X11Y112_SLICE_X14Y112_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B2 = CLBLM_L_X10Y112_SLICE_X13Y112_DQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B3 = CLBLM_L_X10Y107_SLICE_X13Y107_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B4 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D2 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C2 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C3 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C4 = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C5 = CLBLM_R_X11Y110_SLICE_X14Y110_DQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C6 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D3 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D4 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A3 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A4 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_CQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D3 = CLBLM_L_X10Y112_SLICE_X13Y112_DQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D6 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B3 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B4 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A1 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A2 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A3 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A4 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B1 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B2 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B4 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B5 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B6 = CLBLM_L_X8Y112_SLICE_X10Y112_DQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C1 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C2 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C6 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = CLBLL_L_X4Y108_SLICE_X4Y108_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D4 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D1 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_BX = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = CLBLM_R_X7Y107_SLICE_X8Y107_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = CLBLL_L_X4Y108_SLICE_X4Y108_B5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C4 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = CLBLM_R_X5Y108_SLICE_X6Y108_DQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = CLBLL_L_X4Y108_SLICE_X4Y108_DQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A1 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C5 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A4 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_A6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B1 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B2 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B4 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_B6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = CLBLL_L_X4Y108_SLICE_X5Y108_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = CLBLM_R_X5Y112_SLICE_X7Y112_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = CLBLM_R_X5Y108_SLICE_X6Y108_CQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = CLBLL_L_X4Y108_SLICE_X5Y108_CQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = CLBLM_R_X5Y107_SLICE_X7Y107_DQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = CLBLL_L_X4Y108_SLICE_X4Y108_DQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A1 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A2 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A3 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A4 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A5 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A6 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C1 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C2 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_C3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B1 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B2 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B3 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B4 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B5 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B6 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D1 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C2 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C3 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C4 = CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C5 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C6 = CLBLM_R_X7Y106_SLICE_X9Y106_B5Q;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D3 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D4 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X18Y116_D6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D2 = CLBLM_R_X5Y107_SLICE_X7Y107_D5Q;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D3 = CLBLM_R_X11Y107_SLICE_X15Y107_DO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D4 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D5 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B3 = CLBLM_R_X11Y110_SLICE_X15Y110_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B4 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B5 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B6 = CLBLM_R_X11Y110_SLICE_X14Y110_DQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A5 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B1 = CLBLM_R_X11Y112_SLICE_X15Y112_BO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B2 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B6 = CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C1 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C2 = CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C3 = CLBLM_L_X10Y113_SLICE_X12Y113_CQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C5 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D3 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D4 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D5 = CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D3 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D4 = CLBLM_L_X10Y108_SLICE_X12Y108_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A2 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A3 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A6 = CLBLM_L_X8Y109_SLICE_X11Y109_A5Q;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B3 = CLBLM_L_X10Y117_SLICE_X12Y117_DQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B4 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B6 = 1'b1;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C5 = CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C4 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = CLBLL_L_X4Y108_SLICE_X4Y108_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D2 = CLBLM_R_X7Y113_SLICE_X9Y113_DQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D5 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D1 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = CLBLM_R_X3Y110_SLICE_X3Y110_D5Q;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = CLBLM_L_X8Y114_SLICE_X10Y114_D5Q;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C2 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = CLBLM_L_X8Y114_SLICE_X10Y114_D5Q;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A1 = CLBLM_L_X8Y108_SLICE_X11Y108_DQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_AX = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A4 = CLBLM_R_X7Y106_SLICE_X8Y106_DQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = CLBLM_R_X7Y114_SLICE_X8Y114_C5Q;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = CLBLL_L_X4Y109_SLICE_X5Y109_A5Q;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_DQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C1 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C2 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C3 = CLBLM_R_X11Y109_SLICE_X14Y109_A5Q;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = CLBLL_L_X4Y109_SLICE_X5Y109_DQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = CLBLM_R_X5Y107_SLICE_X7Y107_CQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D1 = CLBLM_L_X10Y109_SLICE_X13Y109_BQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D2 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D3 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D4 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D5 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B1 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A1 = CLBLM_L_X10Y107_SLICE_X13Y107_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A2 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A4 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A5 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C1 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C2 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C3 = CLBLM_L_X12Y113_SLICE_X17Y113_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B1 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B2 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B4 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B5 = CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D5 = CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D3 = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C1 = CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C2 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C3 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D4 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C4 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C5 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D3 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D5 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D6 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D1 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D2 = CLBLM_R_X11Y111_SLICE_X15Y111_A5Q;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D3 = CLBLM_R_X11Y107_SLICE_X15Y107_CO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D4 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D5 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D6 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A1 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A3 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A6 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_AX = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B2 = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B5 = CLBLM_L_X10Y113_SLICE_X12Y113_CQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B6 = CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C1 = CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C5 = CLBLM_L_X10Y106_SLICE_X12Y106_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_CO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D3 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D6 = CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A2 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A3 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A6 = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_AX = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B1 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B2 = CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B3 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C2 = CLBLM_L_X10Y114_SLICE_X12Y114_CQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C4 = CLBLM_R_X11Y114_SLICE_X15Y114_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C5 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D1 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D3 = CLBLM_L_X10Y114_SLICE_X12Y114_DQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D5 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = CLBLL_L_X4Y110_SLICE_X5Y110_B5Q;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = CLBLM_R_X5Y107_SLICE_X7Y107_DQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = CLBLL_L_X4Y112_SLICE_X5Y112_BQ;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = CLBLL_L_X4Y108_SLICE_X5Y108_BQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A3 = CLBLM_R_X11Y108_SLICE_X15Y108_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = CLBLL_L_X4Y110_SLICE_X5Y110_CQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = CLBLL_L_X4Y109_SLICE_X5Y109_DQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B2 = CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B3 = CLBLM_L_X12Y108_SLICE_X16Y108_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B4 = CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B6 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = CLBLL_L_X4Y110_SLICE_X5Y110_CQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = CLBLL_L_X4Y109_SLICE_X5Y109_A5Q;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = CLBLL_L_X4Y109_SLICE_X5Y109_DQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C3 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C6 = CLBLM_L_X8Y108_SLICE_X11Y108_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D1 = CLBLM_L_X8Y108_SLICE_X11Y108_CQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D2 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D4 = CLBLM_R_X11Y110_SLICE_X15Y110_BQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D6 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A2 = CLBLM_L_X12Y108_SLICE_X17Y108_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A3 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A6 = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B2 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B4 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B5 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C1 = CLBLM_R_X11Y109_SLICE_X14Y109_A5Q;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C2 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C3 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C5 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C6 = CLBLM_R_X11Y108_SLICE_X14Y108_AQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D1 = CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D2 = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D5 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D6 = CLBLM_R_X11Y109_SLICE_X14Y109_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C4 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C5 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A2 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A3 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A5 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B2 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B5 = CLBLM_L_X12Y114_SLICE_X17Y114_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B6 = CLBLM_L_X10Y110_SLICE_X13Y110_DQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C3 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C4 = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C5 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C6 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D1 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D2 = CLBLM_R_X11Y114_SLICE_X15Y114_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D3 = CLBLM_L_X10Y114_SLICE_X13Y114_DQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D4 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D5 = CLBLM_R_X11Y116_SLICE_X14Y116_DQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D6 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D5 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D6 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A4 = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A6 = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = CLBLM_R_X13Y111_SLICE_X19Y111_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B4 = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_C5Q;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = CLBLM_R_X5Y110_SLICE_X6Y110_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = CLBLM_L_X12Y110_SLICE_X16Y110_D5Q;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_D5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = CLBLM_R_X5Y110_SLICE_X6Y110_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = CLBLL_L_X4Y112_SLICE_X5Y112_C5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D1 = CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D3 = CLBLM_L_X10Y118_SLICE_X12Y118_C5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D5 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = CLBLM_R_X11Y109_SLICE_X14Y109_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A5 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = CLBLL_L_X4Y110_SLICE_X5Y110_CQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A1 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A2 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A3 = CLBLM_L_X10Y107_SLICE_X13Y107_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = CLBLL_L_X4Y111_SLICE_X5Y111_CQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A4 = CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A5 = CLBLM_L_X10Y109_SLICE_X13Y109_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A6 = CLBLM_R_X11Y109_SLICE_X14Y109_BO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B2 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = CLBLM_L_X8Y110_SLICE_X11Y110_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = CLBLL_L_X4Y111_SLICE_X5Y111_DQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C2 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C3 = CLBLM_R_X7Y108_SLICE_X8Y108_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C5 = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C6 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D1 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D2 = CLBLM_L_X8Y108_SLICE_X11Y108_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D4 = CLBLM_L_X12Y112_SLICE_X17Y112_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D5 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A2 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A5 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A6 = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_AX = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B1 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B3 = CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B5 = CLBLM_R_X11Y109_SLICE_X14Y109_A5Q;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C3 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C4 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C5 = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C6 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D1 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D2 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D3 = CLBLM_L_X10Y116_SLICE_X12Y116_DQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D5 = CLBLM_R_X11Y112_SLICE_X14Y112_DQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D6 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C5 = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D4 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D5 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A1 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A3 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A4 = CLBLM_R_X11Y114_SLICE_X15Y114_CQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A6 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_AX = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B1 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B2 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B3 = CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B4 = CLBLM_L_X10Y115_SLICE_X13Y115_CQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B5 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B6 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C2 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C3 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D3 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D4 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A1 = CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A4 = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = CLBLM_R_X11Y109_SLICE_X14Y109_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = CLBLL_L_X4Y108_SLICE_X5Y108_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A3 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A6 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = CLBLM_R_X3Y110_SLICE_X3Y110_CQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B2 = CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B5 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D4 = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D5 = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B6 = CLBLL_L_X4Y108_SLICE_X5Y108_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C4 = CLBLM_R_X7Y106_SLICE_X9Y106_B5Q;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A5 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = CLBLM_R_X5Y109_SLICE_X7Y109_A5Q;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = CLBLL_L_X4Y109_SLICE_X5Y109_A5Q;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = CLBLL_L_X4Y110_SLICE_X5Y110_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = CLBLM_R_X7Y114_SLICE_X8Y114_D5Q;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = CLBLL_L_X4Y109_SLICE_X5Y109_DQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A1 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A3 = CLBLM_R_X11Y110_SLICE_X15Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A4 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A6 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_AX = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B6 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C1 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C5 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D2 = CLBLM_R_X11Y110_SLICE_X15Y110_CQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D3 = CLBLM_L_X10Y107_SLICE_X13Y107_BQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D4 = CLBLM_R_X11Y111_SLICE_X15Y111_A5Q;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D5 = CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A3 = CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A4 = CLBLM_R_X11Y110_SLICE_X15Y110_A5Q;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A5 = CLBLM_R_X11Y110_SLICE_X15Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B1 = CLBLM_L_X12Y113_SLICE_X17Y113_CQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B2 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B3 = CLBLM_R_X11Y109_SLICE_X14Y109_CQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B6 = CLBLM_R_X11Y111_SLICE_X14Y111_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C4 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C5 = CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D1 = CLBLM_R_X11Y110_SLICE_X15Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D2 = CLBLM_R_X11Y110_SLICE_X15Y110_A5Q;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D3 = CLBLM_R_X11Y110_SLICE_X14Y110_DQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D6 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A1 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A2 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A4 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A5 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A1 = CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A2 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A3 = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A6 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = CLBLM_R_X3Y110_SLICE_X3Y110_D5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B1 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B2 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_D5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B4 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B5 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B4 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A1 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A2 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A4 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A5 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_D5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C2 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B1 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B2 = CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B3 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B5 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B6 = CLBLM_R_X7Y107_SLICE_X9Y107_B5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D2 = CLBLM_L_X10Y115_SLICE_X13Y115_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D3 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D4 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D5 = CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D1 = CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C2 = CLBLM_L_X8Y107_SLICE_X11Y107_CQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C3 = CLBLM_L_X8Y107_SLICE_X11Y107_DQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A4 = CLBLM_L_X10Y110_SLICE_X12Y110_DQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A6 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C6 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A1 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A2 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B1 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B2 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B3 = CLBLM_L_X10Y106_SLICE_X12Y106_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B4 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B6 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C2 = CLBLM_L_X8Y117_SLICE_X10Y117_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C4 = CLBLM_R_X13Y116_SLICE_X18Y116_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C6 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A2 = CLBLM_L_X8Y106_SLICE_X10Y106_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = CLBLL_L_X4Y112_SLICE_X4Y112_CQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D2 = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D3 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C2 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C4 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C5 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C6 = CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D1 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D2 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D3 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D4 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D5 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D6 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = CLBLM_L_X10Y113_SLICE_X12Y113_CQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = CLBLL_L_X4Y110_SLICE_X5Y110_CQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = CLBLM_R_X7Y114_SLICE_X9Y114_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A1 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A2 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_C5Q;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A6 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_AX = CLBLM_L_X12Y112_SLICE_X16Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B2 = CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B4 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B6 = CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C2 = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C3 = CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C4 = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C5 = CLBLM_L_X10Y111_SLICE_X12Y111_CQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C6 = CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D2 = CLBLM_L_X10Y111_SLICE_X13Y111_B5Q;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D3 = CLBLM_L_X8Y108_SLICE_X11Y108_DQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D4 = CLBLM_L_X12Y113_SLICE_X16Y113_DQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D6 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_A5Q;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A2 = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A4 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B1 = CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B2 = CLBLM_L_X10Y111_SLICE_X13Y111_DQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B3 = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B4 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B5 = CLBLM_R_X7Y114_SLICE_X8Y114_D5Q;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B6 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C1 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C2 = CLBLM_R_X11Y110_SLICE_X14Y110_CQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C5 = CLBLM_R_X11Y112_SLICE_X15Y112_CQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C6 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_L_X12Y110_SLICE_X16Y110_D5Q;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D1 = CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D2 = CLBLM_L_X10Y111_SLICE_X12Y111_D5Q;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D5 = CLBLM_R_X11Y107_SLICE_X15Y107_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D6 = CLBLM_R_X11Y115_SLICE_X14Y115_DQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_DQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B2 = CLBLM_R_X11Y110_SLICE_X15Y110_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B5 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A1 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A2 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A3 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A4 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A5 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B1 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B3 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B5 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A2 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A3 = CLBLM_L_X8Y108_SLICE_X11Y108_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C4 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C5 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A4 = CLBLM_L_X8Y107_SLICE_X11Y107_CQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A5 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C1 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C2 = CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B2 = CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D3 = CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D4 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D5 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D6 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B6 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D1 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C1 = CLBLM_L_X12Y112_SLICE_X17Y112_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C2 = CLBLM_L_X8Y108_SLICE_X11Y108_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A2 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_C5Q;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A4 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A5 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A6 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B2 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B3 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B4 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B5 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = CLBLL_L_X4Y111_SLICE_X5Y111_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D6 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D6 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C1 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C4 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C5 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A1 = CLBLM_L_X8Y109_SLICE_X10Y109_CQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A4 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B6 = CLBLM_L_X8Y108_SLICE_X11Y108_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C2 = CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C3 = CLBLL_L_X4Y112_SLICE_X5Y112_BQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C6 = CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C5 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D1 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D3 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C6 = CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = CLBLM_L_X10Y114_SLICE_X12Y114_DQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A1 = CLBLM_R_X11Y115_SLICE_X14Y115_CQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A2 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = CLBLM_L_X10Y114_SLICE_X12Y114_DQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B1 = CLBLM_L_X12Y113_SLICE_X17Y113_CQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B2 = CLBLM_L_X12Y110_SLICE_X16Y110_CQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B5 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C2 = CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C5 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C6 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D1 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D2 = CLBLM_L_X12Y112_SLICE_X16Y112_BQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D3 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D4 = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D5 = CLBLM_L_X12Y112_SLICE_X17Y112_BQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D6 = 1'b1;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A1 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A2 = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A3 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A4 = CLBLL_L_X4Y108_SLICE_X5Y108_CQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B2 = CLBLM_R_X11Y112_SLICE_X14Y112_BQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B3 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B4 = CLBLM_R_X11Y110_SLICE_X15Y110_CQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C2 = CLBLM_R_X13Y112_SLICE_X19Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C4 = CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C6 = CLBLM_L_X12Y112_SLICE_X16Y112_A5Q;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D1 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D5 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D6 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A1 = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A2 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A3 = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A6 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B1 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B2 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B3 = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B5 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A1 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A3 = CLBLM_L_X8Y109_SLICE_X11Y109_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A4 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C1 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_AX = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B2 = CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B3 = CLBLM_L_X12Y112_SLICE_X17Y112_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B4 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B6 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D3 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D4 = CLBLM_L_X12Y118_SLICE_X16Y118_AO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D5 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D6 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D1 = CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A1 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A2 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_D5Q;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A4 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A5 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_AX = CLBLM_L_X10Y116_SLICE_X12Y116_D5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_AX = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B1 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B2 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B3 = CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B4 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B5 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_BX = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_D5Q;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C4 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C5 = CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A2 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D1 = CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D5 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B6 = CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C2 = CLBLM_L_X8Y109_SLICE_X10Y109_CQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C4 = CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C5 = CLBLM_R_X7Y114_SLICE_X9Y114_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_SR = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D1 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D2 = CLBLM_L_X8Y111_SLICE_X11Y111_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D5 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = CLBLL_L_X4Y111_SLICE_X5Y111_DQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = CLBLM_R_X5Y108_SLICE_X6Y108_CQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D6 = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = CLBLL_L_X4Y111_SLICE_X5Y111_DQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A1 = CLBLM_L_X8Y108_SLICE_X11Y108_DQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A2 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A3 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B1 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B2 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B4 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_AX = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C1 = CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C2 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C4 = CLBLM_L_X12Y113_SLICE_X16Y113_DQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D2 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D3 = CLBLM_R_X11Y113_SLICE_X15Y113_DQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D6 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A2 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A4 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A5 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A6 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B2 = CLBLM_R_X11Y109_SLICE_X14Y109_CQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B4 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B5 = CLBLM_R_X11Y114_SLICE_X14Y114_BO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C3 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C6 = CLBLM_R_X7Y114_SLICE_X8Y114_DQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D2 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D5 = CLBLM_L_X10Y109_SLICE_X13Y109_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D6 = CLBLM_R_X11Y109_SLICE_X14Y109_CQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A1 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A3 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A5 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A6 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B3 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B4 = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B5 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B6 = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = CLBLM_L_X8Y107_SLICE_X11Y107_CQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = CLBLM_L_X8Y110_SLICE_X11Y110_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C1 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C2 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C3 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = CLBLM_L_X8Y110_SLICE_X11Y110_BQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = CLBLM_L_X8Y109_SLICE_X11Y109_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = CLBLM_L_X8Y109_SLICE_X11Y109_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C2 = CLBLM_L_X8Y106_SLICE_X10Y106_CQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = CLBLM_R_X5Y116_SLICE_X6Y116_A5Q;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = CLBLM_L_X8Y110_SLICE_X11Y110_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = CLBLM_L_X8Y110_SLICE_X11Y110_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_CQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = CLBLL_L_X4Y108_SLICE_X5Y108_CQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A1 = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A2 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A3 = CLBLL_L_X4Y110_SLICE_X5Y110_B5Q;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B1 = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B2 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B6 = CLBLM_L_X10Y114_SLICE_X13Y114_DQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C1 = CLBLM_R_X11Y113_SLICE_X15Y113_CO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C4 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C5 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D1 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D3 = CLBLM_R_X11Y114_SLICE_X15Y114_DQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D4 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A1 = CLBLM_L_X10Y111_SLICE_X13Y111_DQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A4 = CLBLM_L_X10Y114_SLICE_X13Y114_C5Q;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A5 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_AX = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B2 = CLBLM_L_X10Y111_SLICE_X12Y111_D5Q;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B3 = CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C1 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C2 = CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D1 = CLBLM_L_X10Y108_SLICE_X12Y108_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D2 = CLBLM_R_X11Y114_SLICE_X15Y114_DQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D3 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D4 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D5 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_SR = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_A5Q;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = CLBLM_L_X8Y111_SLICE_X11Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = CLBLM_R_X13Y111_SLICE_X18Y111_CQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_DQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = CLBLM_L_X8Y106_SLICE_X10Y106_CQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_C5Q;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = CLBLM_R_X3Y111_SLICE_X3Y111_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A1 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A3 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A4 = CLBLM_L_X12Y116_SLICE_X16Y116_CO5;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A5 = CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A6 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B1 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B2 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B3 = CLBLM_L_X12Y114_SLICE_X16Y114_DQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B4 = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B5 = CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C1 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C2 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C3 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C4 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C5 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D1 = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D2 = CLBLM_R_X13Y115_SLICE_X19Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D3 = CLBLM_R_X11Y116_SLICE_X15Y116_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D4 = CLBLM_R_X11Y115_SLICE_X14Y115_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D5 = CLBLM_R_X13Y115_SLICE_X19Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D6 = CLBLM_R_X13Y116_SLICE_X18Y116_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A2 = CLBLM_L_X10Y115_SLICE_X13Y115_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A3 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A4 = CLBLM_R_X11Y109_SLICE_X14Y109_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B1 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B2 = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B3 = CLBLM_R_X11Y115_SLICE_X14Y115_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C1 = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C3 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C4 = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C6 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D2 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D3 = CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D6 = CLBLM_L_X10Y111_SLICE_X12Y111_D5Q;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B6 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = CLBLM_R_X7Y116_SLICE_X8Y116_C5Q;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A2 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A3 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A5 = CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C1 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_AX = CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C6 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B4 = CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B5 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D3 = CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D5 = CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D6 = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = CLBLM_R_X11Y112_SLICE_X14Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A5 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A6 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C5 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D6 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X4Y112_SLICE_X5Y112_CQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A1 = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A3 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A5 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A6 = CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_AX = CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B1 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B2 = CLBLM_R_X11Y116_SLICE_X15Y116_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B3 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B4 = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B5 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A1 = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A2 = CLBLM_R_X7Y106_SLICE_X9Y106_BQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A5 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C2 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C3 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B2 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_B5Q;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B5 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D1 = CLBLM_L_X12Y116_SLICE_X17Y116_CO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C2 = CLBLM_R_X7Y106_SLICE_X9Y106_CQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C4 = CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C5 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D3 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D4 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A3 = CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A4 = CLBLM_R_X11Y113_SLICE_X15Y113_DQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D3 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D4 = CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D5 = CLBLM_R_X7Y106_SLICE_X9Y106_B5Q;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D6 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B2 = CLBLM_R_X11Y116_SLICE_X14Y116_DQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A3 = CLBLM_R_X7Y106_SLICE_X8Y106_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A6 = CLBLM_R_X7Y106_SLICE_X9Y106_CQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C3 = CLBLM_R_X11Y115_SLICE_X14Y115_B5Q;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B2 = CLBLM_R_X7Y106_SLICE_X8Y106_BQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B3 = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B5 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C2 = CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C3 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C4 = CLBLM_L_X10Y107_SLICE_X13Y107_BQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C6 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D5 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D6 = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B6 = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D2 = CLBLM_R_X7Y106_SLICE_X8Y106_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D3 = CLBLM_R_X7Y106_SLICE_X8Y106_DQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D4 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A3 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A5 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A6 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = CLBLM_L_X12Y114_SLICE_X16Y114_DQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = CLBLM_L_X8Y113_SLICE_X10Y113_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = CLBLM_L_X10Y111_SLICE_X12Y111_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = CLBLM_L_X12Y113_SLICE_X17Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_DQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A2 = CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A4 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A6 = CLBLM_L_X8Y115_SLICE_X11Y115_B5Q;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B2 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B3 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B4 = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B6 = CLBLM_L_X12Y114_SLICE_X17Y114_CQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A1 = CLBLM_L_X8Y108_SLICE_X10Y108_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A2 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A4 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C1 = CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_AX = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C3 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B2 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B4 = CLBLM_R_X7Y109_SLICE_X9Y109_BQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D1 = CLBLM_L_X10Y109_SLICE_X13Y109_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_BX = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D2 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C1 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C3 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C5 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A1 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A2 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A4 = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A5 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D1 = CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D2 = CLBLM_R_X5Y107_SLICE_X7Y107_CQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D4 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D5 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_C5Q;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B1 = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B3 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A2 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A4 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A5 = CLBLM_L_X8Y107_SLICE_X10Y107_DO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A6 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C1 = CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C2 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C3 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B2 = CLBLM_R_X7Y107_SLICE_X8Y107_BQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B4 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D2 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C4 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C5 = CLBLM_R_X5Y107_SLICE_X7Y107_BQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D3 = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D4 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D5 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D6 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D1 = CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D2 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D4 = CLBLM_R_X7Y106_SLICE_X8Y106_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D6 = CLBLM_R_X5Y107_SLICE_X7Y107_BQ;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A3 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A4 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B2 = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B4 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B6 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A2 = CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A6 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B1 = CLBLM_R_X7Y114_SLICE_X8Y114_D5Q;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B6 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C1 = CLBLL_L_X4Y109_SLICE_X5Y109_DQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C2 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C3 = CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D1 = CLBLM_L_X10Y111_SLICE_X12Y111_D5Q;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D2 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D5 = CLBLM_L_X8Y114_SLICE_X10Y114_D5Q;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A1 = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A2 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A3 = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A4 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A5 = CLBLM_L_X8Y109_SLICE_X10Y109_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B1 = CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B2 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B3 = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B5 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B6 = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A1 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A2 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A3 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A4 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C1 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C2 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C3 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B1 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B4 = CLBLM_L_X8Y108_SLICE_X10Y108_AQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B5 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B6 = CLBLM_L_X10Y111_SLICE_X13Y111_DQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C1 = CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C2 = CLBLL_L_X4Y108_SLICE_X4Y108_DQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D1 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C5 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C6 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D2 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A1 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A2 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A3 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A4 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A5 = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D1 = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D2 = CLBLM_R_X7Y106_SLICE_X9Y106_CQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D4 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D4 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D5 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D6 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D5 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_AX = CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B2 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A3 = CLBLM_R_X7Y108_SLICE_X8Y108_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A4 = CLBLM_R_X5Y108_SLICE_X6Y108_BQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C1 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C2 = CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C3 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B1 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B2 = CLBLM_R_X7Y107_SLICE_X8Y107_BQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B3 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D1 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C1 = CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C2 = CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C5 = CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D2 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D3 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D4 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D6 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D1 = CLBLM_L_X8Y108_SLICE_X10Y108_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D4 = CLBLM_L_X10Y111_SLICE_X13Y111_DQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D5 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A3 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A4 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_R_X11Y120_SLICE_X14Y120_A5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B2 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B4 = CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B5 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A1 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A2 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A4 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A5 = CLBLM_R_X3Y111_SLICE_X3Y111_A5Q;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A6 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B2 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B3 = CLBLM_R_X11Y112_SLICE_X14Y112_DQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B4 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C1 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C2 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C3 = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C5 = CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D2 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A1 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A2 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A3 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A5 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_AX = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_C5Q;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B2 = CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B3 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_DQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C4 = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C5 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A4 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C6 = CLBLM_L_X8Y115_SLICE_X10Y115_DO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D1 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D2 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A2 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A3 = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A4 = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A5 = CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B1 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B2 = CLBLM_L_X12Y118_SLICE_X16Y118_AO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B3 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B4 = CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B5 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = CLBLM_L_X8Y111_SLICE_X11Y111_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = CLBLM_L_X8Y113_SLICE_X11Y113_DQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = CLBLM_R_X5Y107_SLICE_X7Y107_CQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B1 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = CLBLM_R_X5Y119_SLICE_X6Y119_A5Q;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C1 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C2 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C3 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = CLBLM_R_X7Y114_SLICE_X8Y114_DQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = CLBLM_R_X5Y112_SLICE_X6Y112_BQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D1 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_DQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D2 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D3 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D4 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D6 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A2 = CLBLM_R_X11Y115_SLICE_X14Y115_B5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A3 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A6 = CLBLM_R_X11Y116_SLICE_X14Y116_C5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_AX = CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B2 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B4 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C1 = CLBLM_R_X11Y115_SLICE_X14Y115_B5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C3 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C4 = CLBLM_R_X11Y116_SLICE_X14Y116_C5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A2 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A5 = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A6 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B1 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B2 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B4 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B5 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B6 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C1 = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C2 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C3 = CLBLM_L_X10Y111_SLICE_X13Y111_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C4 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C5 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A5 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B1 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B3 = CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D1 = CLBLM_R_X11Y116_SLICE_X15Y116_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D2 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D3 = CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D5 = CLBLM_R_X7Y116_SLICE_X8Y116_C5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D3 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = CLBLM_L_X10Y113_SLICE_X12Y113_CQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D5 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A1 = CLBLM_R_X5Y107_SLICE_X7Y107_DQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A2 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A3 = CLBLL_L_X4Y112_SLICE_X5Y112_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A4 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A5 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = CLBLM_R_X5Y117_SLICE_X7Y117_A5Q;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = CLBLM_L_X10Y111_SLICE_X12Y111_BQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = CLBLM_R_X7Y114_SLICE_X8Y114_DQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = CLBLM_R_X7Y106_SLICE_X9Y106_BQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = CLBLM_L_X10Y117_SLICE_X12Y117_DQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A1 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A2 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_D5Q;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A4 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A5 = CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A6 = CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X4Y112_SLICE_X5Y112_C5Q;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C4 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C5 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C6 = CLBLM_L_X10Y115_SLICE_X13Y115_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A2 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A5 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A6 = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_L_X8Y113_SLICE_X10Y113_C5Q;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B1 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B2 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B6 = CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C1 = CLBLM_L_X8Y113_SLICE_X10Y113_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C4 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C5 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D2 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D6 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = CLBLM_L_X12Y112_SLICE_X16Y112_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = CLBLM_R_X7Y114_SLICE_X9Y114_CQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = CLBLM_L_X8Y111_SLICE_X11Y111_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_DQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = CLBLL_L_X4Y108_SLICE_X4Y108_B5Q;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = CLBLM_R_X5Y107_SLICE_X7Y107_DQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = CLBLL_L_X4Y110_SLICE_X5Y110_B5Q;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = CLBLL_L_X4Y112_SLICE_X5Y112_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B1 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B3 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B4 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = CLBLM_L_X8Y115_SLICE_X11Y115_B5Q;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D4 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B6 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D6 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C4 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C2 = CLBLM_R_X11Y114_SLICE_X15Y114_CQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C4 = CLBLM_L_X8Y112_SLICE_X11Y112_BQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C5 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C5 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A1 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A2 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A4 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A5 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C1 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C2 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_D5Q;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C4 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C6 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A4 = CLBLM_L_X10Y111_SLICE_X12Y111_DQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A1 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A2 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A6 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B3 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B1 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B2 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B4 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B6 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = CLBLM_R_X5Y107_SLICE_X7Y107_DQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = CLBLL_L_X4Y112_SLICE_X5Y112_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = CLBLL_L_X4Y110_SLICE_X5Y110_B5Q;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = CLBLL_L_X4Y110_SLICE_X5Y110_B5Q;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C2 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C4 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C5 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = CLBLM_L_X10Y111_SLICE_X12Y111_D5Q;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C6 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = CLBLM_L_X10Y116_SLICE_X12Y116_C5Q;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = CLBLM_L_X8Y115_SLICE_X11Y115_B5Q;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_C5Q;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_AX = CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D3 = CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D6 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D4 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_C5Q;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = CLBLM_R_X7Y114_SLICE_X8Y114_C5Q;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = CLBLM_L_X8Y115_SLICE_X11Y115_B5Q;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A1 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A3 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A5 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A6 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A1 = CLBLM_R_X3Y110_SLICE_X3Y110_DQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A4 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C4 = CLBLM_R_X5Y111_SLICE_X7Y111_CQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = CLBLM_R_X7Y113_SLICE_X9Y113_CQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_AX = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = CLBLM_L_X10Y111_SLICE_X12Y111_D5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = CLBLM_L_X8Y112_SLICE_X11Y112_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_D5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = CLBLM_R_X7Y113_SLICE_X9Y113_DQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = CLBLM_L_X8Y113_SLICE_X10Y113_C5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D3 = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = CLBLM_L_X8Y113_SLICE_X10Y113_DQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_AX = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = CLBLM_L_X8Y113_SLICE_X11Y113_DQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X10Y111_SLICE_X12Y111_DQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = CLBLM_R_X7Y113_SLICE_X8Y113_DQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = CLBLM_R_X11Y112_SLICE_X14Y112_DQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A3 = CLBLM_L_X8Y108_SLICE_X10Y108_AQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B2 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = CLBLM_R_X7Y113_SLICE_X9Y113_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = CLBLM_R_X7Y114_SLICE_X9Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = CLBLM_L_X12Y111_SLICE_X16Y111_B5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = CLBLM_R_X7Y114_SLICE_X9Y114_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = 1'b1;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = CLBLM_L_X10Y111_SLICE_X13Y111_DQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = 1'b1;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B4 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B5 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = CLBLL_L_X4Y108_SLICE_X4Y108_B5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = CLBLM_R_X7Y114_SLICE_X8Y114_DQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = CLBLM_R_X7Y113_SLICE_X8Y113_DQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C5 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D1 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D2 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D3 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A1 = CLBLM_R_X11Y116_SLICE_X14Y116_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A2 = CLBLM_R_X11Y115_SLICE_X14Y115_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A3 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A4 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A1 = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A2 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A4 = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A5 = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B3 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B6 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C2 = CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C3 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C4 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C5 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D2 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D3 = CLBLL_L_X4Y110_SLICE_X5Y110_BQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D5 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A3 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A4 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A5 = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A6 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B1 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B2 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B3 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B4 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B5 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C1 = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C3 = CLBLM_L_X12Y111_SLICE_X16Y111_B5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C4 = CLBLM_R_X13Y115_SLICE_X18Y115_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C6 = CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D2 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D5 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D6 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A3 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A4 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A5 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A6 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B2 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B3 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B4 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B5 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B6 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C3 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C4 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D2 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D3 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D4 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D5 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D6 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B6 = 1'b1;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A6 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A2 = CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A3 = CLBLM_R_X11Y115_SLICE_X14Y115_B5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A5 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A3 = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A5 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B4 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B6 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C3 = CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C4 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D2 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D3 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D4 = CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D5 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A2 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A4 = CLBLM_R_X7Y114_SLICE_X9Y114_C5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A6 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_AX = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B3 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B5 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A1 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A3 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A5 = CLBLM_R_X7Y106_SLICE_X8Y106_BQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A6 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C2 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B2 = CLBLM_R_X5Y107_SLICE_X7Y107_BQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B4 = CLBLL_L_X4Y110_SLICE_X5Y110_BQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B6 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C2 = CLBLM_R_X5Y107_SLICE_X7Y107_CQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C6 = CLBLM_R_X5Y107_SLICE_X7Y107_D5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D3 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D4 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A2 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A3 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A4 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D1 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D4 = CLBLM_R_X7Y107_SLICE_X9Y107_A5Q;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D5 = CLBLL_L_X4Y112_SLICE_X5Y112_BQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B2 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B3 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B4 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B5 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B6 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C2 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_AX = CLBLM_R_X7Y107_SLICE_X8Y107_CO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D2 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D3 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D5 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B4 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B5 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D3 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X4Y112_SLICE_X5Y112_BQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C2 = CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C4 = CLBLM_L_X10Y106_SLICE_X12Y106_BQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A1 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A2 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A3 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A4 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A6 = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B2 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B5 = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B6 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A4 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A5 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A6 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C2 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B2 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B5 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B6 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C1 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C2 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C4 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C6 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D1 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D2 = CLBLM_R_X11Y108_SLICE_X15Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A2 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A3 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A4 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D3 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D5 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D6 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D4 = CLBLM_L_X8Y109_SLICE_X11Y109_A5Q;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D5 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B1 = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B2 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A3 = CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A4 = CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C1 = CLBLM_L_X8Y115_SLICE_X11Y115_B5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C2 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B2 = CLBLM_R_X5Y108_SLICE_X6Y108_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B3 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B6 = CLBLM_R_X3Y114_SLICE_X2Y114_A5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D1 = CLBLM_L_X10Y109_SLICE_X13Y109_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C3 = CLBLM_R_X5Y108_SLICE_X6Y108_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C4 = CLBLM_R_X5Y112_SLICE_X6Y112_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C5 = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D3 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D1 = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D3 = CLBLM_R_X5Y108_SLICE_X6Y108_DQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D4 = CLBLM_R_X13Y109_SLICE_X18Y109_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D5 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D6 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A3 = CLBLM_L_X8Y109_SLICE_X10Y109_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B2 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B3 = CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A5 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B4 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C6 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D1 = CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D3 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D4 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A6 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B6 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = CLBLM_R_X3Y111_SLICE_X3Y111_A5Q;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_AX = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = CLBLM_R_X13Y109_SLICE_X18Y109_CQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = CLBLM_R_X11Y108_SLICE_X14Y108_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = CLBLM_R_X3Y111_SLICE_X3Y111_A5Q;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = CLBLM_R_X5Y112_SLICE_X7Y112_A5Q;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A1 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A2 = CLBLM_L_X8Y117_SLICE_X10Y117_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = CLBLM_L_X8Y113_SLICE_X11Y113_DQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = CLBLM_R_X5Y110_SLICE_X6Y110_BQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A6 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_AX = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B1 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B4 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = CLBLM_R_X11Y107_SLICE_X15Y107_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = CLBLM_R_X11Y108_SLICE_X14Y108_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = CLBLM_R_X7Y114_SLICE_X8Y114_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_L_X12Y110_SLICE_X16Y110_DQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = CLBLL_L_X4Y109_SLICE_X5Y109_A5Q;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = CLBLM_L_X10Y117_SLICE_X12Y117_DQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = CLBLM_R_X7Y109_SLICE_X9Y109_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B5 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C4 = CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C5 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = CLBLM_R_X11Y109_SLICE_X14Y109_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = CLBLM_R_X7Y106_SLICE_X9Y106_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = CLBLL_L_X4Y108_SLICE_X5Y108_BQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D2 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D4 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A4 = CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C3 = CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B4 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B5 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D2 = CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C4 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C4 = CLBLM_R_X13Y115_SLICE_X19Y115_AO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C5 = CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C5 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = CLBLM_R_X7Y109_SLICE_X9Y109_BQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = CLBLM_R_X5Y111_SLICE_X7Y111_CQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = CLBLM_R_X13Y111_SLICE_X18Y111_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = CLBLM_R_X11Y111_SLICE_X14Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = CLBLM_R_X3Y110_SLICE_X3Y110_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = CLBLM_L_X8Y112_SLICE_X11Y112_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y118_SLICE_X17Y118_AQ;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_R_X13Y115_SLICE_X19Y115_AQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B5 = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = CLBLL_L_X4Y111_SLICE_X5Y111_CQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = CLBLM_R_X5Y119_SLICE_X6Y119_A5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = CLBLM_R_X5Y117_SLICE_X7Y117_A5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = CLBLM_R_X7Y114_SLICE_X8Y114_C5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = CLBLM_R_X7Y116_SLICE_X8Y116_C5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_C5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = CLBLM_R_X5Y117_SLICE_X7Y117_A5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = CLBLM_L_X10Y116_SLICE_X12Y116_C5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = CLBLM_R_X5Y119_SLICE_X6Y119_A5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = CLBLM_R_X7Y113_SLICE_X9Y113_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = CLBLM_R_X3Y110_SLICE_X3Y110_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = CLBLM_L_X8Y112_SLICE_X10Y112_DQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = CLBLM_R_X7Y113_SLICE_X9Y113_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = CLBLM_R_X5Y112_SLICE_X6Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = CLBLM_R_X5Y108_SLICE_X6Y108_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_CQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C3 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C6 = CLBLM_L_X8Y109_SLICE_X10Y109_CQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_L_X12Y110_SLICE_X16Y110_D5Q;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D1 = CLBLM_R_X11Y108_SLICE_X15Y108_AQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C4 = CLBLM_R_X11Y116_SLICE_X15Y116_A5Q;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D6 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C4 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = CLBLM_R_X7Y109_SLICE_X9Y109_BQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = CLBLM_R_X7Y113_SLICE_X9Y113_DQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C1 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C2 = CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = CLBLL_L_X4Y109_SLICE_X5Y109_DQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = CLBLM_L_X10Y114_SLICE_X12Y114_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = CLBLM_L_X8Y110_SLICE_X11Y110_AQ;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B5 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A2 = CLBLM_L_X10Y114_SLICE_X13Y114_DQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A4 = CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A5 = CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B2 = CLBLM_R_X5Y109_SLICE_X7Y109_A5Q;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B3 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B4 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B5 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C3 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C6 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A1 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A2 = CLBLM_L_X8Y111_SLICE_X11Y111_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A5 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A6 = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B4 = CLBLM_L_X10Y116_SLICE_X12Y116_C5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B6 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C1 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C2 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C5 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C6 = CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D1 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D3 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D4 = CLBLM_L_X10Y114_SLICE_X13Y114_C5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_L_X12Y110_SLICE_X16Y110_DQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = CLBLL_L_X4Y111_SLICE_X5Y111_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = CLBLM_L_X10Y114_SLICE_X13Y114_DQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = CLBLM_L_X10Y110_SLICE_X13Y110_DQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = CLBLM_R_X5Y111_SLICE_X7Y111_CQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C3 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C4 = CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C5 = CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C6 = CLBLM_L_X12Y114_SLICE_X16Y114_DQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X4Y112_SLICE_X5Y112_CQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = CLBLL_L_X4Y108_SLICE_X5Y108_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D5 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A1 = CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C3 = CLBLM_L_X12Y118_SLICE_X16Y118_AO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C4 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C5 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B3 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D2 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C4 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C5 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X10Y111_SLICE_X12Y111_DQ;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = CLBLM_L_X8Y108_SLICE_X11Y108_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D2 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A3 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D3 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A5 = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D4 = CLBLM_L_X10Y116_SLICE_X12Y116_D5Q;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D6 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C2 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_R_X11Y120_SLICE_X14Y120_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A3 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A4 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B2 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C1 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C2 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C3 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C4 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C5 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C6 = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A1 = CLBLM_R_X5Y119_SLICE_X6Y119_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A2 = CLBLM_R_X5Y116_SLICE_X6Y116_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A3 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A6 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C5 = CLBLM_R_X7Y108_SLICE_X8Y108_AQ;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A4 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B3 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B6 = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C4 = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D3 = CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D4 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D5 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D2 = CLBLM_R_X5Y117_SLICE_X7Y117_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D5 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D6 = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A6 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = CLBLM_L_X8Y111_SLICE_X11Y111_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_AX = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C4 = 1'b1;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X4Y112_SLICE_X5Y112_C5Q;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_L_X8Y113_SLICE_X10Y113_C5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A3 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A4 = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A6 = CLBLL_L_X4Y108_SLICE_X4Y108_DQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B1 = CLBLM_R_X3Y108_SLICE_X2Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B2 = CLBLL_L_X4Y108_SLICE_X4Y108_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B3 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B4 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B5 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B6 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C1 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C2 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C3 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C4 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C5 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C6 = CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A1 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A2 = CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A3 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A4 = CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A5 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D2 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D6 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B2 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B3 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A2 = CLBLM_L_X10Y108_SLICE_X12Y108_BQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A3 = CLBLM_R_X3Y108_SLICE_X2Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A4 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C2 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B2 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B5 = CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B6 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C1 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C2 = CLBLM_R_X3Y108_SLICE_X2Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C3 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C4 = CLBLL_L_X4Y108_SLICE_X4Y108_BQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C5 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D1 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D2 = CLBLM_R_X3Y108_SLICE_X2Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D3 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D4 = CLBLL_L_X4Y108_SLICE_X4Y108_BQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D5 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C4 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C5 = CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C6 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A1 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A3 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_L_X10Y115_SLICE_X12Y115_D5Q;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = CLBLM_R_X5Y108_SLICE_X6Y108_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = CLBLM_L_X10Y109_SLICE_X13Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A1 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A3 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A4 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A6 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_AX = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B1 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B2 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C3 = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D1 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = CLBLM_R_X3Y110_SLICE_X3Y110_D5Q;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = CLBLM_R_X3Y114_SLICE_X2Y114_A5Q;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D3 = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D4 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D5 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = CLBLL_L_X4Y110_SLICE_X4Y110_C5Q;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = CLBLM_R_X3Y110_SLICE_X3Y110_DQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A1 = CLBLM_L_X10Y114_SLICE_X13Y114_A5Q;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C4 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C5 = CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = CLBLM_R_X5Y110_SLICE_X6Y110_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = CLBLL_L_X4Y112_SLICE_X4Y112_DQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C6 = CLBLM_L_X12Y113_SLICE_X17Y113_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B1 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B2 = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C1 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = CLBLM_L_X8Y110_SLICE_X11Y110_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D6 = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = CLBLM_L_X8Y110_SLICE_X11Y110_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D1 = CLBLM_L_X12Y113_SLICE_X17Y113_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D2 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D4 = CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D5 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_SR = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A1 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A2 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X4Y112_SLICE_X5Y112_BQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A3 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A4 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A5 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C4 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B3 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = CLBLM_L_X8Y110_SLICE_X11Y110_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_AX = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = CLBLM_L_X10Y111_SLICE_X12Y111_CQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = CLBLM_R_X7Y106_SLICE_X9Y106_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = CLBLM_R_X3Y111_SLICE_X3Y111_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = CLBLM_R_X3Y110_SLICE_X3Y110_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C1 = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = CLBLM_R_X13Y115_SLICE_X19Y115_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C5 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C6 = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D2 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D5 = CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = CLBLL_L_X4Y109_SLICE_X5Y109_A5Q;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = CLBLM_L_X10Y111_SLICE_X12Y111_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_AX = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D6 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C6 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B5 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B6 = CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D6 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A1 = CLBLM_L_X8Y107_SLICE_X11Y107_DQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A3 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A4 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A6 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D3 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C4 = CLBLM_R_X11Y112_SLICE_X15Y112_CQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B1 = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B4 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B5 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B6 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C5 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C2 = CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C6 = CLBLM_R_X13Y111_SLICE_X19Y111_AQ;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_B6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D4 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D5 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D6 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_C3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_C4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A5 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_C5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = CLBLM_R_X3Y111_SLICE_X3Y111_CQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = CLBLM_R_X11Y115_SLICE_X14Y115_B5Q;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C6 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A4 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B4 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B6 = CLBLM_L_X8Y109_SLICE_X11Y109_A5Q;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_D2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_D3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_CQ;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_D4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_D5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = CLBLM_R_X3Y110_SLICE_X3Y110_DQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C4 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = CLBLM_R_X5Y108_SLICE_X6Y108_DQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A6 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = CLBLM_R_X7Y106_SLICE_X9Y106_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = CLBLL_L_X4Y112_SLICE_X5Y112_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A5 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A1 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A3 = CLBLM_L_X12Y108_SLICE_X17Y108_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A5 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A6 = CLBLM_L_X10Y108_SLICE_X13Y108_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B2 = CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B4 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B5 = CLBLM_L_X12Y108_SLICE_X16Y108_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C6 = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C1 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C2 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C4 = CLBLM_L_X8Y108_SLICE_X11Y108_CQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C6 = CLBLM_R_X13Y109_SLICE_X18Y109_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D1 = CLBLM_L_X10Y108_SLICE_X13Y108_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D2 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D4 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D6 = CLBLM_L_X12Y112_SLICE_X17Y112_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B5 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A1 = CLBLM_R_X11Y108_SLICE_X15Y108_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A3 = CLBLM_L_X12Y108_SLICE_X16Y108_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A6 = CLBLM_R_X11Y109_SLICE_X14Y109_A5Q;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B1 = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B4 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B5 = CLBLM_R_X11Y113_SLICE_X15Y113_DQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B6 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C1 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C3 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C4 = CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = CLBLM_L_X10Y117_SLICE_X12Y117_DQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C5 = CLBLM_R_X11Y110_SLICE_X14Y110_A5Q;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C6 = CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D1 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D2 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D3 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D4 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D5 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D6 = CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C5 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = CLBLM_L_X8Y112_SLICE_X10Y112_DQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y118_SLICE_X17Y118_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_R_X13Y115_SLICE_X19Y115_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A1 = CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A2 = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A4 = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A5 = CLBLM_L_X12Y111_SLICE_X17Y111_CO5;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A6 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B1 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B2 = CLBLM_L_X12Y112_SLICE_X17Y112_AQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B3 = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B4 = CLBLM_L_X10Y108_SLICE_X13Y108_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B5 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B6 = CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C1 = CLBLM_L_X12Y111_SLICE_X17Y111_CO5;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C2 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C4 = CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C5 = CLBLM_R_X13Y109_SLICE_X18Y109_AQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C6 = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLM_R_X37Y115_SLICE_X56Y115_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D1 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D2 = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D3 = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D4 = CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D5 = CLBLM_R_X13Y109_SLICE_X18Y109_AQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A1 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A2 = CLBLM_L_X12Y107_SLICE_X16Y107_DO5;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A3 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A4 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B1 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B2 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B3 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B4 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B5 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C1 = CLBLM_L_X12Y108_SLICE_X17Y108_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C2 = CLBLM_L_X12Y110_SLICE_X16Y110_CQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C3 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C4 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C5 = CLBLM_L_X10Y110_SLICE_X13Y110_CQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C6 = CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D1 = CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D2 = CLBLM_L_X12Y110_SLICE_X16Y110_CQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D3 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D4 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D5 = CLBLM_L_X10Y110_SLICE_X13Y110_CQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C2 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C3 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = CLBLM_R_X5Y112_SLICE_X6Y112_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A3 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A4 = CLBLM_L_X12Y110_SLICE_X17Y110_CQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A5 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A6 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B2 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B4 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B5 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C1 = CLBLM_R_X13Y109_SLICE_X18Y109_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C2 = CLBLM_L_X12Y110_SLICE_X17Y110_CQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C6 = CLBLM_R_X11Y109_SLICE_X14Y109_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D1 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D2 = CLBLM_L_X12Y109_SLICE_X16Y109_BO5;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D3 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D4 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D6 = CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A1 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A3 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A5 = CLBLM_L_X12Y108_SLICE_X17Y108_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A6 = CLBLM_L_X12Y114_SLICE_X16Y114_CQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B2 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B5 = CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B6 = CLBLM_L_X10Y110_SLICE_X13Y110_CQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C1 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C2 = CLBLM_L_X12Y110_SLICE_X16Y110_CQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C4 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D1 = CLBLM_R_X11Y109_SLICE_X14Y109_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D2 = CLBLM_L_X10Y111_SLICE_X13Y111_D5Q;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D3 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D6 = 1'b1;
  assign CLBLM_R_X13Y116_SLICE_X19Y116_D3 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A3 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A4 = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B1 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B4 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B5 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B6 = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C1 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C2 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C3 = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C4 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C6 = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A1 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A4 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A6 = CLBLM_R_X7Y114_SLICE_X9Y114_C5Q;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B1 = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B2 = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B3 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B4 = CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B5 = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B6 = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C5 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C3 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D1 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D3 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A1 = CLBLM_R_X11Y116_SLICE_X15Y116_CQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A2 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A3 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A6 = CLBLM_L_X12Y111_SLICE_X17Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B1 = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B3 = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B4 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B5 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B6 = CLBLM_R_X13Y115_SLICE_X18Y115_BQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C1 = CLBLM_R_X13Y111_SLICE_X19Y111_AQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C2 = CLBLM_R_X13Y111_SLICE_X19Y111_BQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C4 = CLBLM_R_X13Y111_SLICE_X18Y111_BQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C5 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C6 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_A1 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_A2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_A3 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_A4 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_A5 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_A6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D4 = CLBLM_L_X12Y109_SLICE_X16Y109_BO5;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D6 = CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_B1 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_B2 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_B3 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_B4 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_B5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A1 = CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A3 = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A5 = CLBLM_R_X11Y107_SLICE_X15Y107_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A6 = CLBLM_L_X10Y115_SLICE_X12Y115_C5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D3 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_C1 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B1 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B2 = CLBLM_R_X11Y116_SLICE_X15Y116_CQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B3 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B4 = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D6 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X57Y115_D1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C1 = CLBLM_R_X11Y107_SLICE_X15Y107_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C3 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C5 = CLBLM_R_X13Y112_SLICE_X18Y112_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C6 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_A2 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_A3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_A4 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_A6 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_B1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D1 = CLBLM_R_X11Y107_SLICE_X15Y107_BQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D3 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D4 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D5 = CLBLM_L_X12Y113_SLICE_X16Y113_DQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D6 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_B2 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_B3 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_B4 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_B5 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_B6 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_C1 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_C2 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_C3 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_C4 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_C5 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_C6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_D1 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_D2 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_D3 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_D4 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_D5 = 1'b1;
  assign CLBLM_R_X37Y115_SLICE_X56Y115_D6 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C4 = CLBLM_L_X12Y117_SLICE_X16Y117_BO5;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C6 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_AX = CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B2 = 1'b1;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D6 = CLBLM_R_X11Y109_SLICE_X14Y109_CQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A1 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A2 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B2 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B3 = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B4 = CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B5 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B6 = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C1 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C2 = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C3 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C4 = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C5 = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C6 = CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D1 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D2 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D3 = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D4 = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D6 = CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A1 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A3 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A4 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A5 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A6 = CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B4 = CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B6 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C4 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C4 = 1'b1;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D2 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D3 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D4 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D6 = CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A1 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A2 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A3 = CLBLM_L_X12Y112_SLICE_X17Y112_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A5 = CLBLM_L_X12Y110_SLICE_X16Y110_CQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B2 = CLBLM_L_X12Y112_SLICE_X17Y112_BQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B3 = CLBLM_L_X12Y112_SLICE_X16Y112_CO5;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B4 = CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B5 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B6 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B5 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C1 = CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C2 = CLBLM_L_X12Y112_SLICE_X17Y112_CQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C6 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D1 = CLBLM_R_X7Y106_SLICE_X8Y106_DQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D2 = CLBLM_L_X12Y112_SLICE_X17Y112_CQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D3 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D4 = CLBLM_R_X13Y109_SLICE_X18Y109_DQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D5 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A1 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A3 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A4 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A5 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_AX = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B1 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B2 = CLBLM_L_X12Y112_SLICE_X16Y112_BQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B4 = CLBLM_L_X12Y112_SLICE_X16Y112_DO5;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B5 = CLBLM_L_X12Y110_SLICE_X17Y110_CQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B6 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C4 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_BX = CLBLM_L_X12Y112_SLICE_X16Y112_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D5 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C1 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C2 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C4 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C5 = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C5 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C6 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C4 = CLBLM_L_X8Y117_SLICE_X10Y117_CQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D1 = CLBLM_L_X12Y112_SLICE_X17Y112_BQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D2 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D4 = CLBLM_L_X12Y112_SLICE_X16Y112_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D5 = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = CLBLM_L_X10Y117_SLICE_X12Y117_DQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C5 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B5 = CLBLM_R_X7Y119_SLICE_X8Y119_A5Q;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C6 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = CLBLM_L_X10Y114_SLICE_X12Y114_DQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B1 = CLBLM_R_X11Y111_SLICE_X15Y111_A5Q;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B3 = CLBLM_R_X11Y107_SLICE_X15Y107_AQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B4 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A1 = CLBLM_L_X12Y113_SLICE_X17Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A2 = CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A3 = CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A5 = CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A6 = CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B3 = CLBLM_R_X13Y112_SLICE_X18Y112_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B5 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C1 = CLBLM_R_X13Y118_SLICE_X18Y118_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C2 = CLBLM_L_X12Y113_SLICE_X17Y113_CQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C5 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C4 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D1 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D3 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D5 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C5 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A1 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A2 = CLBLM_L_X12Y114_SLICE_X16Y114_BQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A3 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A5 = CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A6 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B1 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B2 = CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B4 = CLBLM_R_X7Y113_SLICE_X8Y113_DQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C2 = CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C4 = CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C5 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C6 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D5 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D6 = 1'b1;
endmodule
