module top(
  input LIOB33_SING_X0Y0_IOB_X0Y0_IPAD,
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_SING_X0Y149_IOB_X0Y149_IPAD,
  input LIOB33_SING_X0Y150_IOB_X0Y150_IPAD,
  input LIOB33_SING_X0Y199_IOB_X0Y199_IPAD,
  input LIOB33_SING_X0Y200_IOB_X0Y200_IPAD,
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_SING_X0Y99_IOB_X0Y99_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y119_IOB_X0Y119_IPAD,
  input LIOB33_X0Y119_IOB_X0Y120_IPAD,
  input LIOB33_X0Y11_IOB_X0Y11_IPAD,
  input LIOB33_X0Y11_IOB_X0Y12_IPAD,
  input LIOB33_X0Y121_IOB_X0Y121_IPAD,
  input LIOB33_X0Y121_IOB_X0Y122_IPAD,
  input LIOB33_X0Y123_IOB_X0Y123_IPAD,
  input LIOB33_X0Y123_IOB_X0Y124_IPAD,
  input LIOB33_X0Y125_IOB_X0Y125_IPAD,
  input LIOB33_X0Y125_IOB_X0Y126_IPAD,
  input LIOB33_X0Y127_IOB_X0Y127_IPAD,
  input LIOB33_X0Y127_IOB_X0Y128_IPAD,
  input LIOB33_X0Y129_IOB_X0Y129_IPAD,
  input LIOB33_X0Y129_IOB_X0Y130_IPAD,
  input LIOB33_X0Y131_IOB_X0Y131_IPAD,
  input LIOB33_X0Y131_IOB_X0Y132_IPAD,
  input LIOB33_X0Y133_IOB_X0Y133_IPAD,
  input LIOB33_X0Y133_IOB_X0Y134_IPAD,
  input LIOB33_X0Y135_IOB_X0Y135_IPAD,
  input LIOB33_X0Y135_IOB_X0Y136_IPAD,
  input LIOB33_X0Y137_IOB_X0Y137_IPAD,
  input LIOB33_X0Y137_IOB_X0Y138_IPAD,
  input LIOB33_X0Y139_IOB_X0Y139_IPAD,
  input LIOB33_X0Y139_IOB_X0Y140_IPAD,
  input LIOB33_X0Y13_IOB_X0Y13_IPAD,
  input LIOB33_X0Y13_IOB_X0Y14_IPAD,
  input LIOB33_X0Y141_IOB_X0Y141_IPAD,
  input LIOB33_X0Y141_IOB_X0Y142_IPAD,
  input LIOB33_X0Y143_IOB_X0Y143_IPAD,
  input LIOB33_X0Y145_IOB_X0Y145_IPAD,
  input LIOB33_X0Y145_IOB_X0Y146_IPAD,
  input LIOB33_X0Y147_IOB_X0Y147_IPAD,
  input LIOB33_X0Y147_IOB_X0Y148_IPAD,
  input LIOB33_X0Y151_IOB_X0Y151_IPAD,
  input LIOB33_X0Y151_IOB_X0Y152_IPAD,
  input LIOB33_X0Y153_IOB_X0Y153_IPAD,
  input LIOB33_X0Y153_IOB_X0Y154_IPAD,
  input LIOB33_X0Y155_IOB_X0Y155_IPAD,
  input LIOB33_X0Y155_IOB_X0Y156_IPAD,
  input LIOB33_X0Y157_IOB_X0Y157_IPAD,
  input LIOB33_X0Y157_IOB_X0Y158_IPAD,
  input LIOB33_X0Y159_IOB_X0Y159_IPAD,
  input LIOB33_X0Y159_IOB_X0Y160_IPAD,
  input LIOB33_X0Y15_IOB_X0Y15_IPAD,
  input LIOB33_X0Y15_IOB_X0Y16_IPAD,
  input LIOB33_X0Y161_IOB_X0Y161_IPAD,
  input LIOB33_X0Y161_IOB_X0Y162_IPAD,
  input LIOB33_X0Y163_IOB_X0Y163_IPAD,
  input LIOB33_X0Y163_IOB_X0Y164_IPAD,
  input LIOB33_X0Y165_IOB_X0Y165_IPAD,
  input LIOB33_X0Y165_IOB_X0Y166_IPAD,
  input LIOB33_X0Y167_IOB_X0Y167_IPAD,
  input LIOB33_X0Y167_IOB_X0Y168_IPAD,
  input LIOB33_X0Y169_IOB_X0Y169_IPAD,
  input LIOB33_X0Y169_IOB_X0Y170_IPAD,
  input LIOB33_X0Y171_IOB_X0Y171_IPAD,
  input LIOB33_X0Y171_IOB_X0Y172_IPAD,
  input LIOB33_X0Y173_IOB_X0Y173_IPAD,
  input LIOB33_X0Y173_IOB_X0Y174_IPAD,
  input LIOB33_X0Y175_IOB_X0Y175_IPAD,
  input LIOB33_X0Y175_IOB_X0Y176_IPAD,
  input LIOB33_X0Y177_IOB_X0Y177_IPAD,
  input LIOB33_X0Y177_IOB_X0Y178_IPAD,
  input LIOB33_X0Y179_IOB_X0Y179_IPAD,
  input LIOB33_X0Y179_IOB_X0Y180_IPAD,
  input LIOB33_X0Y17_IOB_X0Y17_IPAD,
  input LIOB33_X0Y17_IOB_X0Y18_IPAD,
  input LIOB33_X0Y181_IOB_X0Y181_IPAD,
  input LIOB33_X0Y181_IOB_X0Y182_IPAD,
  input LIOB33_X0Y183_IOB_X0Y183_IPAD,
  input LIOB33_X0Y183_IOB_X0Y184_IPAD,
  input LIOB33_X0Y185_IOB_X0Y185_IPAD,
  input LIOB33_X0Y185_IOB_X0Y186_IPAD,
  input LIOB33_X0Y187_IOB_X0Y187_IPAD,
  input LIOB33_X0Y187_IOB_X0Y188_IPAD,
  input LIOB33_X0Y189_IOB_X0Y189_IPAD,
  input LIOB33_X0Y189_IOB_X0Y190_IPAD,
  input LIOB33_X0Y191_IOB_X0Y191_IPAD,
  input LIOB33_X0Y191_IOB_X0Y192_IPAD,
  input LIOB33_X0Y193_IOB_X0Y193_IPAD,
  input LIOB33_X0Y193_IOB_X0Y194_IPAD,
  input LIOB33_X0Y195_IOB_X0Y195_IPAD,
  input LIOB33_X0Y195_IOB_X0Y196_IPAD,
  input LIOB33_X0Y197_IOB_X0Y197_IPAD,
  input LIOB33_X0Y197_IOB_X0Y198_IPAD,
  input LIOB33_X0Y19_IOB_X0Y19_IPAD,
  input LIOB33_X0Y19_IOB_X0Y20_IPAD,
  input LIOB33_X0Y1_IOB_X0Y1_IPAD,
  input LIOB33_X0Y1_IOB_X0Y2_IPAD,
  input LIOB33_X0Y201_IOB_X0Y201_IPAD,
  input LIOB33_X0Y201_IOB_X0Y202_IPAD,
  input LIOB33_X0Y203_IOB_X0Y203_IPAD,
  input LIOB33_X0Y203_IOB_X0Y204_IPAD,
  input LIOB33_X0Y205_IOB_X0Y205_IPAD,
  input LIOB33_X0Y205_IOB_X0Y206_IPAD,
  input LIOB33_X0Y207_IOB_X0Y207_IPAD,
  input LIOB33_X0Y207_IOB_X0Y208_IPAD,
  input LIOB33_X0Y209_IOB_X0Y209_IPAD,
  input LIOB33_X0Y209_IOB_X0Y210_IPAD,
  input LIOB33_X0Y211_IOB_X0Y211_IPAD,
  input LIOB33_X0Y211_IOB_X0Y212_IPAD,
  input LIOB33_X0Y213_IOB_X0Y213_IPAD,
  input LIOB33_X0Y213_IOB_X0Y214_IPAD,
  input LIOB33_X0Y215_IOB_X0Y215_IPAD,
  input LIOB33_X0Y215_IOB_X0Y216_IPAD,
  input LIOB33_X0Y217_IOB_X0Y217_IPAD,
  input LIOB33_X0Y217_IOB_X0Y218_IPAD,
  input LIOB33_X0Y219_IOB_X0Y219_IPAD,
  input LIOB33_X0Y219_IOB_X0Y220_IPAD,
  input LIOB33_X0Y21_IOB_X0Y21_IPAD,
  input LIOB33_X0Y21_IOB_X0Y22_IPAD,
  input LIOB33_X0Y221_IOB_X0Y221_IPAD,
  input LIOB33_X0Y221_IOB_X0Y222_IPAD,
  input LIOB33_X0Y223_IOB_X0Y223_IPAD,
  input LIOB33_X0Y223_IOB_X0Y224_IPAD,
  input LIOB33_X0Y225_IOB_X0Y225_IPAD,
  input LIOB33_X0Y225_IOB_X0Y226_IPAD,
  input LIOB33_X0Y227_IOB_X0Y227_IPAD,
  input LIOB33_X0Y227_IOB_X0Y228_IPAD,
  input LIOB33_X0Y229_IOB_X0Y229_IPAD,
  input LIOB33_X0Y229_IOB_X0Y230_IPAD,
  input LIOB33_X0Y231_IOB_X0Y231_IPAD,
  input LIOB33_X0Y231_IOB_X0Y232_IPAD,
  input LIOB33_X0Y233_IOB_X0Y233_IPAD,
  input LIOB33_X0Y233_IOB_X0Y234_IPAD,
  input LIOB33_X0Y235_IOB_X0Y235_IPAD,
  input LIOB33_X0Y235_IOB_X0Y236_IPAD,
  input LIOB33_X0Y237_IOB_X0Y237_IPAD,
  input LIOB33_X0Y237_IOB_X0Y238_IPAD,
  input LIOB33_X0Y239_IOB_X0Y239_IPAD,
  input LIOB33_X0Y239_IOB_X0Y240_IPAD,
  input LIOB33_X0Y23_IOB_X0Y23_IPAD,
  input LIOB33_X0Y23_IOB_X0Y24_IPAD,
  input LIOB33_X0Y241_IOB_X0Y241_IPAD,
  input LIOB33_X0Y241_IOB_X0Y242_IPAD,
  input LIOB33_X0Y243_IOB_X0Y243_IPAD,
  input LIOB33_X0Y25_IOB_X0Y25_IPAD,
  input LIOB33_X0Y25_IOB_X0Y26_IPAD,
  input LIOB33_X0Y27_IOB_X0Y27_IPAD,
  input LIOB33_X0Y27_IOB_X0Y28_IPAD,
  input LIOB33_X0Y3_IOB_X0Y3_IPAD,
  input LIOB33_X0Y3_IOB_X0Y4_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y5_IOB_X0Y5_IPAD,
  input LIOB33_X0Y5_IOB_X0Y6_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input LIOB33_X0Y79_IOB_X0Y80_IPAD,
  input LIOB33_X0Y7_IOB_X0Y7_IPAD,
  input LIOB33_X0Y7_IOB_X0Y8_IPAD,
  input LIOB33_X0Y81_IOB_X0Y81_IPAD,
  input LIOB33_X0Y81_IOB_X0Y82_IPAD,
  input LIOB33_X0Y83_IOB_X0Y83_IPAD,
  input LIOB33_X0Y83_IOB_X0Y84_IPAD,
  input LIOB33_X0Y85_IOB_X0Y85_IPAD,
  input LIOB33_X0Y85_IOB_X0Y86_IPAD,
  input LIOB33_X0Y87_IOB_X0Y87_IPAD,
  input LIOB33_X0Y87_IOB_X0Y88_IPAD,
  input LIOB33_X0Y89_IOB_X0Y89_IPAD,
  input LIOB33_X0Y89_IOB_X0Y90_IPAD,
  input LIOB33_X0Y91_IOB_X0Y91_IPAD,
  input LIOB33_X0Y91_IOB_X0Y92_IPAD,
  input LIOB33_X0Y93_IOB_X0Y93_IPAD,
  input LIOB33_X0Y93_IOB_X0Y94_IPAD,
  input LIOB33_X0Y95_IOB_X0Y95_IPAD,
  input LIOB33_X0Y95_IOB_X0Y96_IPAD,
  input LIOB33_X0Y97_IOB_X0Y97_IPAD,
  input LIOB33_X0Y97_IOB_X0Y98_IPAD,
  input LIOB33_X0Y9_IOB_X0Y10_IPAD,
  input LIOB33_X0Y9_IOB_X0Y9_IPAD,
  input RIOB33_SING_X105Y150_IOB_X1Y150_IPAD,
  input RIOB33_X105Y151_IOB_X1Y151_IPAD,
  input RIOB33_X105Y151_IOB_X1Y152_IPAD,
  input RIOB33_X105Y153_IOB_X1Y153_IPAD,
  input RIOB33_X105Y153_IOB_X1Y154_IPAD,
  input RIOB33_X105Y155_IOB_X1Y155_IPAD,
  input RIOB33_X105Y155_IOB_X1Y156_IPAD,
  input RIOB33_X105Y157_IOB_X1Y157_IPAD,
  input RIOB33_X105Y157_IOB_X1Y158_IPAD,
  input RIOB33_X105Y159_IOB_X1Y159_IPAD,
  output RIOB33_SING_X105Y100_IOB_X1Y100_OPAD,
  output RIOB33_SING_X105Y149_IOB_X1Y149_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_SING_X105Y50_IOB_X1Y50_OPAD,
  output RIOB33_SING_X105Y99_IOB_X1Y99_OPAD,
  output RIOB33_X105Y101_IOB_X1Y101_OPAD,
  output RIOB33_X105Y101_IOB_X1Y102_OPAD,
  output RIOB33_X105Y103_IOB_X1Y103_OPAD,
  output RIOB33_X105Y103_IOB_X1Y104_OPAD,
  output RIOB33_X105Y105_IOB_X1Y105_OPAD,
  output RIOB33_X105Y105_IOB_X1Y106_OPAD,
  output RIOB33_X105Y107_IOB_X1Y107_OPAD,
  output RIOB33_X105Y107_IOB_X1Y108_OPAD,
  output RIOB33_X105Y109_IOB_X1Y109_OPAD,
  output RIOB33_X105Y109_IOB_X1Y110_OPAD,
  output RIOB33_X105Y111_IOB_X1Y111_OPAD,
  output RIOB33_X105Y111_IOB_X1Y112_OPAD,
  output RIOB33_X105Y113_IOB_X1Y113_OPAD,
  output RIOB33_X105Y113_IOB_X1Y114_OPAD,
  output RIOB33_X105Y115_IOB_X1Y115_OPAD,
  output RIOB33_X105Y115_IOB_X1Y116_OPAD,
  output RIOB33_X105Y117_IOB_X1Y117_OPAD,
  output RIOB33_X105Y117_IOB_X1Y118_OPAD,
  output RIOB33_X105Y119_IOB_X1Y119_OPAD,
  output RIOB33_X105Y119_IOB_X1Y120_OPAD,
  output RIOB33_X105Y121_IOB_X1Y121_OPAD,
  output RIOB33_X105Y121_IOB_X1Y122_OPAD,
  output RIOB33_X105Y123_IOB_X1Y123_OPAD,
  output RIOB33_X105Y123_IOB_X1Y124_OPAD,
  output RIOB33_X105Y125_IOB_X1Y125_OPAD,
  output RIOB33_X105Y125_IOB_X1Y126_OPAD,
  output RIOB33_X105Y127_IOB_X1Y127_OPAD,
  output RIOB33_X105Y127_IOB_X1Y128_OPAD,
  output RIOB33_X105Y129_IOB_X1Y129_OPAD,
  output RIOB33_X105Y129_IOB_X1Y130_OPAD,
  output RIOB33_X105Y131_IOB_X1Y131_OPAD,
  output RIOB33_X105Y131_IOB_X1Y132_OPAD,
  output RIOB33_X105Y133_IOB_X1Y133_OPAD,
  output RIOB33_X105Y133_IOB_X1Y134_OPAD,
  output RIOB33_X105Y135_IOB_X1Y135_OPAD,
  output RIOB33_X105Y135_IOB_X1Y136_OPAD,
  output RIOB33_X105Y137_IOB_X1Y137_OPAD,
  output RIOB33_X105Y137_IOB_X1Y138_OPAD,
  output RIOB33_X105Y139_IOB_X1Y139_OPAD,
  output RIOB33_X105Y139_IOB_X1Y140_OPAD,
  output RIOB33_X105Y141_IOB_X1Y141_OPAD,
  output RIOB33_X105Y141_IOB_X1Y142_OPAD,
  output RIOB33_X105Y143_IOB_X1Y143_OPAD,
  output RIOB33_X105Y143_IOB_X1Y144_OPAD,
  output RIOB33_X105Y145_IOB_X1Y145_OPAD,
  output RIOB33_X105Y145_IOB_X1Y146_OPAD,
  output RIOB33_X105Y147_IOB_X1Y147_OPAD,
  output RIOB33_X105Y147_IOB_X1Y148_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD,
  output RIOB33_X105Y51_IOB_X1Y51_OPAD,
  output RIOB33_X105Y51_IOB_X1Y52_OPAD,
  output RIOB33_X105Y53_IOB_X1Y53_OPAD,
  output RIOB33_X105Y53_IOB_X1Y54_OPAD,
  output RIOB33_X105Y55_IOB_X1Y55_OPAD,
  output RIOB33_X105Y55_IOB_X1Y56_OPAD,
  output RIOB33_X105Y57_IOB_X1Y57_OPAD,
  output RIOB33_X105Y57_IOB_X1Y58_OPAD,
  output RIOB33_X105Y59_IOB_X1Y59_OPAD,
  output RIOB33_X105Y59_IOB_X1Y60_OPAD,
  output RIOB33_X105Y61_IOB_X1Y61_OPAD,
  output RIOB33_X105Y61_IOB_X1Y62_OPAD,
  output RIOB33_X105Y63_IOB_X1Y63_OPAD,
  output RIOB33_X105Y63_IOB_X1Y64_OPAD,
  output RIOB33_X105Y65_IOB_X1Y65_OPAD,
  output RIOB33_X105Y65_IOB_X1Y66_OPAD,
  output RIOB33_X105Y67_IOB_X1Y67_OPAD,
  output RIOB33_X105Y67_IOB_X1Y68_OPAD,
  output RIOB33_X105Y69_IOB_X1Y69_OPAD,
  output RIOB33_X105Y69_IOB_X1Y70_OPAD,
  output RIOB33_X105Y71_IOB_X1Y71_OPAD,
  output RIOB33_X105Y71_IOB_X1Y72_OPAD,
  output RIOB33_X105Y73_IOB_X1Y73_OPAD,
  output RIOB33_X105Y73_IOB_X1Y74_OPAD,
  output RIOB33_X105Y75_IOB_X1Y75_OPAD,
  output RIOB33_X105Y75_IOB_X1Y76_OPAD,
  output RIOB33_X105Y77_IOB_X1Y77_OPAD,
  output RIOB33_X105Y77_IOB_X1Y78_OPAD,
  output RIOB33_X105Y79_IOB_X1Y79_OPAD,
  output RIOB33_X105Y79_IOB_X1Y80_OPAD,
  output RIOB33_X105Y81_IOB_X1Y81_OPAD,
  output RIOB33_X105Y81_IOB_X1Y82_OPAD,
  output RIOB33_X105Y83_IOB_X1Y83_OPAD,
  output RIOB33_X105Y83_IOB_X1Y84_OPAD,
  output RIOB33_X105Y85_IOB_X1Y85_OPAD,
  output RIOB33_X105Y85_IOB_X1Y86_OPAD,
  output RIOB33_X105Y87_IOB_X1Y87_OPAD,
  output RIOB33_X105Y87_IOB_X1Y88_OPAD,
  output RIOB33_X105Y89_IOB_X1Y89_OPAD,
  output RIOB33_X105Y89_IOB_X1Y90_OPAD,
  output RIOB33_X105Y91_IOB_X1Y91_OPAD,
  output RIOB33_X105Y91_IOB_X1Y92_OPAD,
  output RIOB33_X105Y93_IOB_X1Y93_OPAD,
  output RIOB33_X105Y93_IOB_X1Y94_OPAD,
  output RIOB33_X105Y95_IOB_X1Y95_OPAD,
  output RIOB33_X105Y95_IOB_X1Y96_OPAD,
  output RIOB33_X105Y97_IOB_X1Y97_OPAD,
  output RIOB33_X105Y97_IOB_X1Y98_OPAD
  );
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_AO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_AO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_BO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_CO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_CO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_DO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_DO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_AO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_BO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_BO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_CO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_CO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_DO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_DO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_AO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_BO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_CO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_DO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_AO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_BO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_DO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_BO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_CO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_DO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_AO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_BO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_DO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_DO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_AO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_AO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_BO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_BO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_CO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_DO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_DO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_AO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_BO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_BO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_CO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_CO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_DO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_DO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_AO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_AO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_BO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_BO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_CO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_CO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_DO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_DO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_DO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_DO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_BO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_BO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_DO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_DO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_AO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_AO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_BO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_BO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_DO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_DO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_DO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_AMUX;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_AO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_AO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_BO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_BO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_CO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_CO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_DO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_DO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AMUX;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_BMUX;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_BO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_CO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_CO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_DO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_DO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_AO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_BO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_BO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_CO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_DO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_DO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_BO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_BO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_DO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_DO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_AO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_AO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_BO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_DO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_DO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_AO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_BO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_CO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_CO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_DO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_DO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_AO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_AO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_BO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_BO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_CO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_CO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_DO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_DO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_CO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_DO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_DO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D_XOR;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_A;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_A1;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_A2;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_A3;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_A4;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_A5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_A6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_AO5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_AO6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_A_CY;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_A_XOR;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_B;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_B1;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_B2;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_B3;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_B4;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_B5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_B6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_BO5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_BO6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_B_CY;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_B_XOR;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_C;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_C1;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_C2;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_C3;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_C4;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_C5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_C6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_CO5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_CO6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_C_CY;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_C_XOR;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_D;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_D1;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_D2;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_D3;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_D4;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_D5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_D6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_DO5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_DO6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_D_CY;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X0Y165_D_XOR;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_A;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_A1;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_A2;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_A3;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_A4;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_A5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_A6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_AO5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_AO6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_A_CY;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_A_XOR;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_B;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_B1;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_B2;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_B3;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_B4;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_B5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_B6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_BO5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_BO6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_B_CY;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_B_XOR;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_C;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_C1;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_C2;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_C3;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_C4;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_C5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_C6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_CO5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_CO6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_C_CY;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_C_XOR;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_D;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_D1;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_D2;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_D3;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_D4;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_D5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_D6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_DO5;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_DO6;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_D_CY;
  wire [0:0] CLBLL_L_X2Y165_SLICE_X1Y165_D_XOR;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_A;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_A1;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_A2;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_A3;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_A4;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_A5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_A6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_AO5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_AO6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_A_CY;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_A_XOR;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_B;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_B1;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_B2;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_B3;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_B4;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_B5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_B6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_BO5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_BO6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_B_CY;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_B_XOR;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_C;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_C1;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_C2;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_C3;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_C4;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_C5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_C6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_CO5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_CO6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_C_CY;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_C_XOR;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_D;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_D1;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_D2;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_D3;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_D4;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_D5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_D6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_DO5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_DO6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_D_CY;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X0Y170_D_XOR;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_A;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_A1;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_A2;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_A3;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_A4;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_A5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_A6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_AO5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_AO6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_A_CY;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_A_XOR;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_B;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_B1;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_B2;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_B3;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_B4;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_B5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_B6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_BO5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_BO6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_B_CY;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_B_XOR;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_C;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_C1;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_C2;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_C3;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_C4;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_C5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_C6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_CO5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_CO6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_C_CY;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_C_XOR;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_D;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_D1;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_D2;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_D3;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_D4;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_D5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_D6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_DO5;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_DO6;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_D_CY;
  wire [0:0] CLBLL_L_X2Y170_SLICE_X1Y170_D_XOR;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_A;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_A1;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_A2;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_A3;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_A4;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_A5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_A6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_AMUX;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_AO5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_AO6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_A_CY;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_A_XOR;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_B;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_B1;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_B2;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_B3;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_B4;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_B5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_B6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_BO5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_BO6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_B_CY;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_B_XOR;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_C;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_C1;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_C2;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_C3;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_C4;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_C5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_C6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_CO5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_CO6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_C_CY;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_C_XOR;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_D;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_D1;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_D2;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_D3;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_D4;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_D5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_D6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_DO5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_DO6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_D_CY;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X0Y187_D_XOR;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_A;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_A1;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_A2;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_A3;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_A4;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_A5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_A6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_AO5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_AO6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_A_CY;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_A_XOR;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_B;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_B1;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_B2;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_B3;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_B4;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_B5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_B6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_BO5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_BO6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_B_CY;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_B_XOR;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_C;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_C1;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_C2;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_C3;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_C4;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_C5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_C6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_CO5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_CO6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_C_CY;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_C_XOR;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_D;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_D1;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_D2;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_D3;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_D4;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_D5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_D6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_DO5;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_DO6;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_D_CY;
  wire [0:0] CLBLL_L_X2Y187_SLICE_X1Y187_D_XOR;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_A;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_A1;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_A2;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_A3;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_A4;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_A5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_A6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_AO5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_AO6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_A_CY;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_A_XOR;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_B;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_B1;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_B2;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_B3;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_B4;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_B5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_B6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_BO5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_BO6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_B_CY;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_B_XOR;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_C;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_C1;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_C2;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_C3;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_C4;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_C5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_C6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_CO5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_CO6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_C_CY;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_C_XOR;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_D;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_D1;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_D2;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_D3;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_D4;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_D5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_D6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_DO5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_DO6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_D_CY;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X0Y189_D_XOR;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_A;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_A1;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_A2;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_A3;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_A4;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_A5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_A6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_AO5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_AO6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_A_CY;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_A_XOR;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_B;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_B1;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_B2;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_B3;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_B4;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_B5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_B6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_BO5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_BO6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_B_CY;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_B_XOR;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_C;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_C1;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_C2;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_C3;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_C4;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_C5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_C6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_CO5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_CO6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_C_CY;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_C_XOR;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_D;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_D1;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_D2;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_D3;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_D4;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_D5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_D6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_DO5;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_DO6;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_D_CY;
  wire [0:0] CLBLL_L_X2Y189_SLICE_X1Y189_D_XOR;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_A;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_A1;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_A2;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_A3;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_A4;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_A5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_A6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_AO5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_AO6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_A_CY;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_A_XOR;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_B;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_B1;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_B2;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_B3;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_B4;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_B5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_B6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_BO5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_BO6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_B_CY;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_B_XOR;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_C;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_C1;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_C2;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_C3;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_C4;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_C5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_C6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_CO5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_CO6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_C_CY;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_C_XOR;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_D;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_D1;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_D2;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_D3;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_D4;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_D5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_D6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_DO5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_DO6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_D_CY;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X0Y192_D_XOR;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_A;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_A1;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_A2;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_A3;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_A4;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_A5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_A6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_AO5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_AO6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_A_CY;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_A_XOR;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_B;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_B1;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_B2;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_B3;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_B4;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_B5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_B6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_BO5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_BO6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_B_CY;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_B_XOR;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_C;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_C1;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_C2;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_C3;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_C4;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_C5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_C6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_CO5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_CO6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_C_CY;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_C_XOR;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_D;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_D1;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_D2;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_D3;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_D4;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_D5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_D6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_DO5;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_DO6;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_D_CY;
  wire [0:0] CLBLL_L_X2Y192_SLICE_X1Y192_D_XOR;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_A;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_A1;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_A2;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_A3;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_A4;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_A5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_A6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_AO5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_AO6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_A_CY;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_A_XOR;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_B;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_B1;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_B2;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_B3;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_B4;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_B5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_B6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_BO5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_BO6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_B_CY;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_B_XOR;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_C;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_C1;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_C2;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_C3;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_C4;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_C5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_C6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_CO5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_CO6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_C_CY;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_C_XOR;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_D;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_D1;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_D2;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_D3;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_D4;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_D5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_D6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_DO5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_DO6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_D_CY;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X0Y193_D_XOR;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_A;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_A1;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_A2;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_A3;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_A4;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_A5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_A6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_AO5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_AO6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_A_CY;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_A_XOR;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_B;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_B1;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_B2;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_B3;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_B4;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_B5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_B6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_BO5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_BO6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_B_CY;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_B_XOR;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_C;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_C1;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_C2;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_C3;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_C4;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_C5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_C6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_CO5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_CO6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_C_CY;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_C_XOR;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_D;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_D1;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_D2;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_D3;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_D4;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_D5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_D6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_DO5;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_DO6;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_D_CY;
  wire [0:0] CLBLL_L_X2Y193_SLICE_X1Y193_D_XOR;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_A;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_A1;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_A2;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_A3;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_A4;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_A5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_A6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_AO5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_AO6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_A_CY;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_A_XOR;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_B;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_B1;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_B2;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_B3;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_B4;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_B5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_B6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_BO5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_BO6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_B_CY;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_B_XOR;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_C;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_C1;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_C2;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_C3;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_C4;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_C5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_C6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_CO5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_CO6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_C_CY;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_C_XOR;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_D;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_D1;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_D2;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_D3;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_D4;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_D5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_D6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_DO5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_DO6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_D_CY;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X0Y194_D_XOR;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_A;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_A1;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_A2;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_A3;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_A4;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_A5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_A6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_AO5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_AO6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_A_CY;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_A_XOR;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_B;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_B1;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_B2;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_B3;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_B4;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_B5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_B6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_BO5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_BO6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_B_CY;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_B_XOR;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_C;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_C1;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_C2;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_C3;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_C4;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_C5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_C6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_CO5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_CO6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_C_CY;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_C_XOR;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_D;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_D1;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_D2;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_D3;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_D4;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_D5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_D6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_DO5;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_DO6;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_D_CY;
  wire [0:0] CLBLL_L_X2Y194_SLICE_X1Y194_D_XOR;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_A;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_A1;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_A2;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_A3;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_A4;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_A5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_A6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_AO5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_AO6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_A_CY;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_A_XOR;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_B;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_B1;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_B2;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_B3;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_B4;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_B5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_B6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_BO5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_BO6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_B_CY;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_B_XOR;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_C;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_C1;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_C2;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_C3;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_C4;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_C5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_C6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_CO5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_CO6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_C_CY;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_C_XOR;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_D;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_D1;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_D2;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_D3;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_D4;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_D5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_D6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_DO5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_DO6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_D_CY;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X0Y208_D_XOR;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_A;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_A1;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_A2;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_A3;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_A4;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_A5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_A6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_AO5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_AO6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_A_CY;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_A_XOR;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_B;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_B1;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_B2;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_B3;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_B4;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_B5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_B6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_BO5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_BO6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_B_CY;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_B_XOR;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_C;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_C1;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_C2;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_C3;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_C4;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_C5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_C6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_CO5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_CO6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_C_CY;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_C_XOR;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_D;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_D1;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_D2;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_D3;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_D4;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_D5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_D6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_DO5;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_DO6;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_D_CY;
  wire [0:0] CLBLL_L_X2Y208_SLICE_X1Y208_D_XOR;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_A;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_A1;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_A2;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_A3;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_A4;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_A5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_A6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_AO5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_AO6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_A_CY;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_A_XOR;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_B;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_B1;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_B2;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_B3;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_B4;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_B5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_B6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_BO5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_BO6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_B_CY;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_B_XOR;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_C;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_C1;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_C2;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_C3;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_C4;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_C5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_C6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_CO5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_CO6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_C_CY;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_C_XOR;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_D;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_D1;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_D2;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_D3;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_D4;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_D5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_D6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_DO5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_DO6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_D_CY;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X0Y210_D_XOR;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_A;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_A1;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_A2;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_A3;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_A4;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_A5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_A6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_AO5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_AO6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_A_CY;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_A_XOR;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_B;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_B1;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_B2;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_B3;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_B4;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_B5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_B6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_BO5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_BO6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_B_CY;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_B_XOR;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_C;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_C1;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_C2;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_C3;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_C4;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_C5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_C6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_CO5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_CO6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_C_CY;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_C_XOR;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_D;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_D1;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_D2;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_D3;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_D4;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_D5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_D6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_DO5;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_DO6;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_D_CY;
  wire [0:0] CLBLL_L_X2Y210_SLICE_X1Y210_D_XOR;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_A;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_A1;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_A2;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_A3;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_A4;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_A5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_A6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_AMUX;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_AO5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_AO6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_A_CY;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_A_XOR;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_B;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_B1;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_B2;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_B3;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_B4;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_B5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_B6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_BO5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_BO6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_B_CY;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_B_XOR;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_C;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_C1;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_C2;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_C3;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_C4;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_C5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_C6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_CO5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_CO6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_C_CY;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_C_XOR;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_D;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_D1;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_D2;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_D3;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_D4;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_D5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_D6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_DO5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_DO6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_D_CY;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X66Y152_D_XOR;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_A;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_A1;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_A2;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_A3;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_A4;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_A5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_A6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_AO5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_AO6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_A_CY;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_A_XOR;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_B;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_B1;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_B2;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_B3;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_B4;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_B5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_B6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_BO5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_BO6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_B_CY;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_B_XOR;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_C;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_C1;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_C2;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_C3;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_C4;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_C5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_C6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_CO5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_CO6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_C_CY;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_C_XOR;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_D;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_D1;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_D2;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_D3;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_D4;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_D5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_D6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_DO5;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_DO6;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_D_CY;
  wire [0:0] CLBLM_L_X44Y152_SLICE_X67Y152_D_XOR;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_A;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_A1;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_A2;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_A3;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_A4;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_A5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_A6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_AMUX;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_AO5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_AO6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_A_CY;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_A_XOR;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_B;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_B1;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_B2;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_B3;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_B4;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_B5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_B6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_BMUX;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_BO5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_BO6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_B_CY;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_B_XOR;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_C;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_C1;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_C2;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_C3;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_C4;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_C5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_C6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_CO5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_CO6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_C_CY;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_C_XOR;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_D;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_D1;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_D2;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_D3;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_D4;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_D5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_D6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_DO5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_DO6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_D_CY;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X66Y158_D_XOR;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_A;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_A1;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_A2;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_A3;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_A4;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_A5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_A6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_AO5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_AO6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_A_CY;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_A_XOR;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_B;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_B1;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_B2;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_B3;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_B4;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_B5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_B6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_BO5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_BO6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_B_CY;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_B_XOR;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_C;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_C1;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_C2;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_C3;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_C4;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_C5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_C6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_CO5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_CO6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_C_CY;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_C_XOR;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_D;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_D1;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_D2;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_D3;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_D4;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_D5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_D6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_DO5;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_DO6;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_D_CY;
  wire [0:0] CLBLM_L_X44Y158_SLICE_X67Y158_D_XOR;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_A;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_A1;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_A2;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_A3;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_A4;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_A5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_A6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_AO5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_AO6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_A_CY;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_A_XOR;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_B;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_B1;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_B2;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_B3;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_B4;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_B5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_B6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_BO5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_BO6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_B_CY;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_B_XOR;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_C;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_C1;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_C2;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_C3;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_C4;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_C5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_C6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_CO5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_CO6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_C_CY;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_C_XOR;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_D;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_D1;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_D2;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_D3;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_D4;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_D5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_D6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_DO5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_DO6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_D_CY;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X72Y145_D_XOR;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_A;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_A1;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_A2;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_A3;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_A4;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_A5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_A6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_AO5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_AO6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_A_CY;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_A_XOR;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_B;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_B1;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_B2;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_B3;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_B4;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_B5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_B6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_BO5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_BO6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_B_CY;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_B_XOR;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_C;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_C1;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_C2;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_C3;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_C4;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_C5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_C6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_CO5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_CO6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_C_CY;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_C_XOR;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_D;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_D1;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_D2;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_D3;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_D4;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_D5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_D6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_DO5;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_DO6;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_D_CY;
  wire [0:0] CLBLM_R_X47Y145_SLICE_X73Y145_D_XOR;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_A;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_A1;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_A2;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_A3;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_A4;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_A5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_A6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_AMUX;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_AO5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_AO6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_A_CY;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_A_XOR;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_B;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_B1;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_B2;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_B3;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_B4;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_B5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_B6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_BO5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_BO6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_B_CY;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_B_XOR;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_C;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_C1;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_C2;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_C3;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_C4;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_C5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_C6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_CO5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_CO6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_C_CY;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_C_XOR;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_D;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_D1;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_D2;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_D3;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_D4;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_D5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_D6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_DO5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_DO6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_D_CY;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X72Y158_D_XOR;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_A;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_A1;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_A2;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_A3;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_A4;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_A5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_A6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_AO5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_AO6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_A_CY;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_A_XOR;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_B;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_B1;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_B2;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_B3;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_B4;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_B5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_B6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_BO5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_BO6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_B_CY;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_B_XOR;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_C;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_C1;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_C2;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_C3;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_C4;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_C5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_C6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_CO5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_CO6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_C_CY;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_C_XOR;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_D;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_D1;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_D2;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_D3;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_D4;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_D5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_D6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_DO5;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_DO6;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_D_CY;
  wire [0:0] CLBLM_R_X47Y158_SLICE_X73Y158_D_XOR;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_A;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_A1;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_A2;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_A3;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_A4;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_A5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_A6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_AO5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_AO6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_A_CY;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_A_XOR;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_B;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_B1;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_B2;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_B3;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_B4;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_B5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_B6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_BO5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_BO6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_B_CY;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_B_XOR;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_C;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_C1;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_C2;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_C3;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_C4;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_C5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_C6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_CO5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_CO6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_C_CY;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_C_XOR;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_D;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_D1;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_D2;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_D3;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_D4;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_D5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_D6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_DO5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_DO6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_D_CY;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X88Y133_D_XOR;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_A;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_A1;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_A2;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_A3;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_A4;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_A5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_A6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_AO5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_AO6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_A_CY;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_A_XOR;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_B;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_B1;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_B2;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_B3;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_B4;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_B5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_B6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_BO5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_BO6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_B_CY;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_B_XOR;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_C;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_C1;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_C2;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_C3;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_C4;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_C5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_C6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_CO5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_CO6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_C_CY;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_C_XOR;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_D;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_D1;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_D2;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_D3;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_D4;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_D5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_D6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_DO5;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_DO6;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_D_CY;
  wire [0:0] CLBLM_R_X59Y133_SLICE_X89Y133_D_XOR;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_A;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_A1;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_A2;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_A3;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_A4;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_A5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_A6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_AO5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_AO6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_A_CY;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_A_XOR;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_B;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_B1;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_B2;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_B3;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_B4;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_B5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_B6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_BO5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_BO6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_B_CY;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_B_XOR;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_C;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_C1;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_C2;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_C3;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_C4;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_C5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_C6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_CO5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_CO6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_C_CY;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_C_XOR;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_D;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_D1;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_D2;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_D3;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_D4;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_D5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_D6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_DO5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_DO6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_D_CY;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X88Y159_D_XOR;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_A;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_A1;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_A2;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_A3;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_A4;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_A5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_A6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_AO5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_AO6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_A_CY;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_A_XOR;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_B;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_B1;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_B2;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_B3;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_B4;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_B5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_B6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_BO5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_BO6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_B_CY;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_B_XOR;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_C;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_C1;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_C2;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_C3;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_C4;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_C5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_C6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_CO5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_CO6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_C_CY;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_C_XOR;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_D;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_D1;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_D2;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_D3;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_D4;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_D5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_D6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_DO5;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_DO6;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_D_CY;
  wire [0:0] CLBLM_R_X59Y159_SLICE_X89Y159_D_XOR;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_A;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_A1;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_A2;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_A3;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_A4;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_A5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_A6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_AO5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_AO6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_A_CY;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_A_XOR;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_B;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_B1;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_B2;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_B3;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_B4;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_B5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_B6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_BO5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_BO6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_B_CY;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_B_XOR;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_C;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_C1;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_C2;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_C3;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_C4;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_C5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_C6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_CO5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_CO6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_C_CY;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_C_XOR;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_D;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_D1;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_D2;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_D3;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_D4;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_D5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_D6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_DO5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_DO6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_D_CY;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X100Y130_D_XOR;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_A;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_A1;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_A2;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_A3;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_A4;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_A5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_A6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_AO5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_AO6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_A_CY;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_A_XOR;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_B;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_B1;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_B2;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_B3;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_B4;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_B5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_B6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_BO5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_BO6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_B_CY;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_B_XOR;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_C;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_C1;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_C2;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_C3;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_C4;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_C5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_C6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_CO5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_CO6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_C_CY;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_C_XOR;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_D;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_D1;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_D2;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_D3;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_D4;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_D5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_D6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_DO5;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_DO6;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_D_CY;
  wire [0:0] CLBLM_R_X67Y130_SLICE_X101Y130_D_XOR;
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_I;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_I;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_I;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_I;
  wire [0:0] LIOB33_SING_X0Y200_IOB_X0Y200_I;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_SING_X0Y99_IOB_X0Y99_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y12_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_I;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_I;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_I;
  wire [0:0] LIOB33_X0Y13_IOB_X0Y13_I;
  wire [0:0] LIOB33_X0Y13_IOB_X0Y14_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_I;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_I;
  wire [0:0] LIOB33_X0Y15_IOB_X0Y15_I;
  wire [0:0] LIOB33_X0Y15_IOB_X0Y16_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_I;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_I;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y17_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y18_I;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_I;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_I;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_I;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_I;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_I;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_I;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_I;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_I;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_I;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_I;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_I;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_I;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_I;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_I;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_I;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_I;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_I;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_I;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y19_I;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y20_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_I;
  wire [0:0] LIOB33_X0Y201_IOB_X0Y201_I;
  wire [0:0] LIOB33_X0Y201_IOB_X0Y202_I;
  wire [0:0] LIOB33_X0Y203_IOB_X0Y203_I;
  wire [0:0] LIOB33_X0Y203_IOB_X0Y204_I;
  wire [0:0] LIOB33_X0Y205_IOB_X0Y205_I;
  wire [0:0] LIOB33_X0Y205_IOB_X0Y206_I;
  wire [0:0] LIOB33_X0Y207_IOB_X0Y207_I;
  wire [0:0] LIOB33_X0Y207_IOB_X0Y208_I;
  wire [0:0] LIOB33_X0Y209_IOB_X0Y209_I;
  wire [0:0] LIOB33_X0Y209_IOB_X0Y210_I;
  wire [0:0] LIOB33_X0Y211_IOB_X0Y211_I;
  wire [0:0] LIOB33_X0Y211_IOB_X0Y212_I;
  wire [0:0] LIOB33_X0Y213_IOB_X0Y213_I;
  wire [0:0] LIOB33_X0Y213_IOB_X0Y214_I;
  wire [0:0] LIOB33_X0Y215_IOB_X0Y215_I;
  wire [0:0] LIOB33_X0Y215_IOB_X0Y216_I;
  wire [0:0] LIOB33_X0Y217_IOB_X0Y217_I;
  wire [0:0] LIOB33_X0Y217_IOB_X0Y218_I;
  wire [0:0] LIOB33_X0Y219_IOB_X0Y219_I;
  wire [0:0] LIOB33_X0Y219_IOB_X0Y220_I;
  wire [0:0] LIOB33_X0Y21_IOB_X0Y21_I;
  wire [0:0] LIOB33_X0Y21_IOB_X0Y22_I;
  wire [0:0] LIOB33_X0Y221_IOB_X0Y221_I;
  wire [0:0] LIOB33_X0Y221_IOB_X0Y222_I;
  wire [0:0] LIOB33_X0Y223_IOB_X0Y223_I;
  wire [0:0] LIOB33_X0Y223_IOB_X0Y224_I;
  wire [0:0] LIOB33_X0Y225_IOB_X0Y225_I;
  wire [0:0] LIOB33_X0Y225_IOB_X0Y226_I;
  wire [0:0] LIOB33_X0Y227_IOB_X0Y227_I;
  wire [0:0] LIOB33_X0Y227_IOB_X0Y228_I;
  wire [0:0] LIOB33_X0Y229_IOB_X0Y229_I;
  wire [0:0] LIOB33_X0Y229_IOB_X0Y230_I;
  wire [0:0] LIOB33_X0Y231_IOB_X0Y231_I;
  wire [0:0] LIOB33_X0Y231_IOB_X0Y232_I;
  wire [0:0] LIOB33_X0Y233_IOB_X0Y233_I;
  wire [0:0] LIOB33_X0Y233_IOB_X0Y234_I;
  wire [0:0] LIOB33_X0Y235_IOB_X0Y235_I;
  wire [0:0] LIOB33_X0Y235_IOB_X0Y236_I;
  wire [0:0] LIOB33_X0Y237_IOB_X0Y237_I;
  wire [0:0] LIOB33_X0Y237_IOB_X0Y238_I;
  wire [0:0] LIOB33_X0Y239_IOB_X0Y239_I;
  wire [0:0] LIOB33_X0Y239_IOB_X0Y240_I;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y23_I;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y24_I;
  wire [0:0] LIOB33_X0Y241_IOB_X0Y241_I;
  wire [0:0] LIOB33_X0Y241_IOB_X0Y242_I;
  wire [0:0] LIOB33_X0Y243_IOB_X0Y243_I;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y25_I;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y26_I;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y27_I;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y28_I;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_I;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y4_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y5_I;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y6_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y7_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y8_I;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y81_I;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y82_I;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y83_I;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y84_I;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y85_I;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y86_I;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y87_I;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y88_I;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y89_I;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y90_I;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y91_I;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y92_I;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y93_I;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y94_I;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y95_I;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y96_I;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y97_I;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y98_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y10_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y9_I;
  wire [0:0] LIOI3_SING_X0Y0_ILOGIC_X0Y0_D;
  wire [0:0] LIOI3_SING_X0Y0_ILOGIC_X0Y0_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_ILOGIC_X0Y149_D;
  wire [0:0] LIOI3_SING_X0Y149_ILOGIC_X0Y149_O;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_D;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_O;
  wire [0:0] LIOI3_SING_X0Y199_ILOGIC_X0Y199_D;
  wire [0:0] LIOI3_SING_X0Y199_ILOGIC_X0Y199_O;
  wire [0:0] LIOI3_SING_X0Y200_ILOGIC_X0Y200_D;
  wire [0:0] LIOI3_SING_X0Y200_ILOGIC_X0Y200_O;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_SING_X0Y99_ILOGIC_X0Y99_D;
  wire [0:0] LIOI3_SING_X0Y99_ILOGIC_X0Y99_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y207_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y207_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y208_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y208_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y219_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y219_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y220_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y220_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y231_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y231_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y232_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y232_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y243_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y243_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y213_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y213_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y214_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y214_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y237_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y237_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y238_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y238_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y136_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y136_O;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y139_D;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y139_O;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y140_D;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y140_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_O;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y148_D;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y148_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_O;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_D;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_O;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_D;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_O;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y168_D;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y168_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y178_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y178_O;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y179_D;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y179_O;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y180_D;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y180_O;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_D;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_O;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_D;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_O;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y183_D;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y183_O;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y184_D;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y184_O;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y185_D;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y185_O;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y186_D;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y186_O;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y189_D;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y189_O;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y190_D;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y190_O;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y191_D;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y191_O;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y192_D;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y192_O;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y195_D;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y195_O;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y196_D;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y196_O;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y197_D;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y197_O;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y198_D;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y198_O;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y1_D;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y1_O;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y2_D;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y2_O;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y201_D;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y201_O;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y202_D;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y202_O;
  wire [0:0] LIOI3_X0Y203_ILOGIC_X0Y203_D;
  wire [0:0] LIOI3_X0Y203_ILOGIC_X0Y203_O;
  wire [0:0] LIOI3_X0Y203_ILOGIC_X0Y204_D;
  wire [0:0] LIOI3_X0Y203_ILOGIC_X0Y204_O;
  wire [0:0] LIOI3_X0Y205_ILOGIC_X0Y205_D;
  wire [0:0] LIOI3_X0Y205_ILOGIC_X0Y205_O;
  wire [0:0] LIOI3_X0Y205_ILOGIC_X0Y206_D;
  wire [0:0] LIOI3_X0Y205_ILOGIC_X0Y206_O;
  wire [0:0] LIOI3_X0Y209_ILOGIC_X0Y209_D;
  wire [0:0] LIOI3_X0Y209_ILOGIC_X0Y209_O;
  wire [0:0] LIOI3_X0Y209_ILOGIC_X0Y210_D;
  wire [0:0] LIOI3_X0Y209_ILOGIC_X0Y210_O;
  wire [0:0] LIOI3_X0Y211_ILOGIC_X0Y211_D;
  wire [0:0] LIOI3_X0Y211_ILOGIC_X0Y211_O;
  wire [0:0] LIOI3_X0Y211_ILOGIC_X0Y212_D;
  wire [0:0] LIOI3_X0Y211_ILOGIC_X0Y212_O;
  wire [0:0] LIOI3_X0Y215_ILOGIC_X0Y215_D;
  wire [0:0] LIOI3_X0Y215_ILOGIC_X0Y215_O;
  wire [0:0] LIOI3_X0Y215_ILOGIC_X0Y216_D;
  wire [0:0] LIOI3_X0Y215_ILOGIC_X0Y216_O;
  wire [0:0] LIOI3_X0Y217_ILOGIC_X0Y217_D;
  wire [0:0] LIOI3_X0Y217_ILOGIC_X0Y217_O;
  wire [0:0] LIOI3_X0Y217_ILOGIC_X0Y218_D;
  wire [0:0] LIOI3_X0Y217_ILOGIC_X0Y218_O;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_D;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_O;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_D;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_O;
  wire [0:0] LIOI3_X0Y221_ILOGIC_X0Y222_D;
  wire [0:0] LIOI3_X0Y221_ILOGIC_X0Y222_O;
  wire [0:0] LIOI3_X0Y223_ILOGIC_X0Y223_D;
  wire [0:0] LIOI3_X0Y223_ILOGIC_X0Y223_O;
  wire [0:0] LIOI3_X0Y223_ILOGIC_X0Y224_D;
  wire [0:0] LIOI3_X0Y223_ILOGIC_X0Y224_O;
  wire [0:0] LIOI3_X0Y225_ILOGIC_X0Y225_D;
  wire [0:0] LIOI3_X0Y225_ILOGIC_X0Y225_O;
  wire [0:0] LIOI3_X0Y225_ILOGIC_X0Y226_D;
  wire [0:0] LIOI3_X0Y225_ILOGIC_X0Y226_O;
  wire [0:0] LIOI3_X0Y227_ILOGIC_X0Y227_D;
  wire [0:0] LIOI3_X0Y227_ILOGIC_X0Y227_O;
  wire [0:0] LIOI3_X0Y227_ILOGIC_X0Y228_D;
  wire [0:0] LIOI3_X0Y227_ILOGIC_X0Y228_O;
  wire [0:0] LIOI3_X0Y229_ILOGIC_X0Y229_D;
  wire [0:0] LIOI3_X0Y229_ILOGIC_X0Y229_O;
  wire [0:0] LIOI3_X0Y229_ILOGIC_X0Y230_D;
  wire [0:0] LIOI3_X0Y229_ILOGIC_X0Y230_O;
  wire [0:0] LIOI3_X0Y233_ILOGIC_X0Y234_D;
  wire [0:0] LIOI3_X0Y233_ILOGIC_X0Y234_O;
  wire [0:0] LIOI3_X0Y235_ILOGIC_X0Y235_D;
  wire [0:0] LIOI3_X0Y235_ILOGIC_X0Y235_O;
  wire [0:0] LIOI3_X0Y235_ILOGIC_X0Y236_D;
  wire [0:0] LIOI3_X0Y235_ILOGIC_X0Y236_O;
  wire [0:0] LIOI3_X0Y239_ILOGIC_X0Y239_D;
  wire [0:0] LIOI3_X0Y239_ILOGIC_X0Y239_O;
  wire [0:0] LIOI3_X0Y239_ILOGIC_X0Y240_D;
  wire [0:0] LIOI3_X0Y239_ILOGIC_X0Y240_O;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_D;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_O;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_D;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_O;
  wire [0:0] LIOI3_X0Y241_ILOGIC_X0Y241_D;
  wire [0:0] LIOI3_X0Y241_ILOGIC_X0Y241_O;
  wire [0:0] LIOI3_X0Y241_ILOGIC_X0Y242_D;
  wire [0:0] LIOI3_X0Y241_ILOGIC_X0Y242_O;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_D;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_O;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_D;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_O;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_D;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_O;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_D;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_O;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y3_D;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y3_O;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y4_D;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y4_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_O;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y80_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y80_O;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y83_D;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y83_O;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y84_D;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y84_O;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y85_D;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y85_O;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y86_D;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y86_O;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y89_D;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y89_O;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y90_D;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y90_O;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y91_D;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y91_O;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y92_D;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y92_O;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y95_D;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y95_O;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y96_D;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y96_O;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y97_D;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y97_O;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y98_D;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y98_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_O;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_O;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_I;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_SING_X105Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_SING_X105Y99_IOB_X1Y99_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_I;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_I;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_I;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_I;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_I;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_I;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_I;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_I;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y53_O;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y54_O;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y56_O;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y57_O;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y59_O;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y60_O;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y62_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y63_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y64_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y65_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y66_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y67_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y68_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y69_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y70_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y71_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y72_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y73_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y74_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y75_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y76_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y77_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y78_O;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y79_O;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y80_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y81_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y82_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y83_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y84_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y85_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y86_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y87_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y88_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y89_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y90_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y91_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y92_O;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y93_O;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y94_O;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y95_O;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y96_O;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y97_O;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y98_O;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ;
  wire [0:0] RIOI3_SING_X105Y150_ILOGIC_X1Y150_D;
  wire [0:0] RIOI3_SING_X105Y150_ILOGIC_X1Y150_O;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_D1;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_OQ;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_T1;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_TQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_TQ;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y151_D;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y151_O;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y152_D;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y152_O;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y153_D;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y153_O;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y154_D;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y154_O;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y155_D;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y155_O;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y156_D;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y156_O;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y159_D;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y159_O;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_D1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_OQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_T1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_TQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_D1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_OQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_T1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_TQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_D1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_OQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_T1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_TQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_D1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_OQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_T1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_TQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_D1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_OQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_T1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_TQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_D1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_OQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_T1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_TQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_D1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_OQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_T1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_TQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_D1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_OQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_T1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_TQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_D1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_OQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_T1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_TQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_D1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_OQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_T1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_TQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_D1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_OQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_T1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_TQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_D1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_OQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_T1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_DO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_CO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_BO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfc)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y13_IOB_X0Y14_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(1'b1),
.I4(RIOB33_X105Y155_IOB_X1Y156_I),
.I5(LIOB33_X0Y5_IOB_X0Y5_I),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_AO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_DO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_CO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_BO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_AO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000110011)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(LIOB33_X0Y51_IOB_X0Y51_I),
.I2(1'b1),
.I3(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.I4(1'b1),
.I5(RIOB33_X105Y155_IOB_X1Y155_I),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_DO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000100010001)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y153_IOB_X1Y154_I),
.I2(LIOB33_X0Y3_IOB_X0Y4_I),
.I3(LIOB33_X0Y13_IOB_X0Y13_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_CO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00ff01)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_BLUT (
.I0(LIOB33_X0Y17_IOB_X0Y17_I),
.I1(RIOB33_X105Y157_IOB_X1Y158_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y163_IOB_X0Y164_I),
.I4(LIOB33_X0Y7_IOB_X0Y7_I),
.I5(LIOB33_X0Y161_IOB_X0Y162_I),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_BO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccffccffcd)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_ALUT (
.I0(LIOB33_X0Y51_IOB_X0Y51_I),
.I1(LIOB33_X0Y163_IOB_X0Y164_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y161_IOB_X0Y162_I),
.I4(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.I5(RIOB33_X105Y155_IOB_X1Y155_I),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_AO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_DO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_CO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033333332)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_BLUT (
.I0(LIOB33_X0Y3_IOB_X0Y4_I),
.I1(LIOB33_X0Y161_IOB_X0Y162_I),
.I2(LIOB33_X0Y13_IOB_X0Y13_I),
.I3(RIOB33_X105Y153_IOB_X1Y154_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(LIOB33_X0Y163_IOB_X0Y164_I),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_BO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccffccffcd)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_ALUT (
.I0(LIOB33_X0Y3_IOB_X0Y4_I),
.I1(LIOB33_X0Y161_IOB_X0Y162_I),
.I2(LIOB33_X0Y13_IOB_X0Y13_I),
.I3(LIOB33_X0Y163_IOB_X0Y164_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y153_IOB_X1Y154_I),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_AO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_DO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000100010001)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_CLUT (
.I0(LIOB33_X0Y151_IOB_X0Y151_I),
.I1(LIOB33_X0Y11_IOB_X0Y12_I),
.I2(LIOB33_X0Y3_IOB_X0Y3_I),
.I3(RIOB33_X105Y153_IOB_X1Y153_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_CO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010115055)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_BLUT (
.I0(CLBLL_L_X2Y103_SLICE_X0Y103_DO6),
.I1(CLBLL_L_X2Y103_SLICE_X0Y103_CO6),
.I2(CLBLL_L_X2Y102_SLICE_X0Y102_AO6),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I4(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I5(CLBLL_L_X2Y104_SLICE_X0Y104_CO6),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_BO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0fff0fff1)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_ALUT (
.I0(LIOB33_X0Y11_IOB_X0Y12_I),
.I1(LIOB33_X0Y3_IOB_X0Y3_I),
.I2(LIOB33_X0Y161_IOB_X0Y162_I),
.I3(LIOB33_X0Y163_IOB_X0Y164_I),
.I4(LIOB33_X0Y151_IOB_X0Y151_I),
.I5(RIOB33_X105Y153_IOB_X1Y153_I),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_AO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_DO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_CO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_BO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_AO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000505)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_ALUT (
.I0(LIOB33_X0Y1_IOB_X0Y2_I),
.I1(1'b1),
.I2(LIOB33_X0Y243_IOB_X0Y243_I),
.I3(1'b1),
.I4(LIOB33_X0Y11_IOB_X0Y11_I),
.I5(RIOB33_X105Y151_IOB_X1Y152_I),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_DO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000000f)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_SING_X0Y0_IOB_X0Y0_I),
.I3(RIOB33_X105Y151_IOB_X1Y151_I),
.I4(LIOB33_X0Y241_IOB_X0Y241_I),
.I5(LIOB33_X0Y9_IOB_X0Y9_I),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_BO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0fff0fff1)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_ALUT (
.I0(LIOB33_X0Y9_IOB_X0Y9_I),
.I1(LIOB33_SING_X0Y0_IOB_X0Y0_I),
.I2(LIOB33_X0Y161_IOB_X0Y162_I),
.I3(LIOB33_X0Y163_IOB_X0Y164_I),
.I4(LIOB33_X0Y241_IOB_X0Y241_I),
.I5(RIOB33_X105Y151_IOB_X1Y151_I),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_AO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_DO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_CO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_BO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_AO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff0f)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(1'b1),
.I4(LIOB33_X0Y131_IOB_X0Y131_I),
.I5(LIOB33_X0Y123_IOB_X0Y124_I),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_DO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000011)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_CLUT (
.I0(LIOB33_X0Y151_IOB_X0Y152_I),
.I1(RIOB33_X105Y157_IOB_X1Y157_I),
.I2(1'b1),
.I3(LIOB33_X0Y5_IOB_X0Y6_I),
.I4(LIOB33_X0Y15_IOB_X0Y16_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_CO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033333332)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_BLUT (
.I0(LIOB33_X0Y17_IOB_X0Y18_I),
.I1(CLBLL_L_X2Y103_SLICE_X0Y103_BO6),
.I2(RIOB33_SING_X105Y150_IOB_X1Y150_I),
.I3(LIOB33_X0Y7_IOB_X0Y8_I),
.I4(RIOB33_X105Y159_IOB_X1Y159_I),
.I5(LIOB33_X0Y179_IOB_X0Y180_I),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_BO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff00fe00)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_ALUT (
.I0(CLBLL_L_X2Y104_SLICE_X0Y104_BO6),
.I1(LIOB33_X0Y15_IOB_X0Y16_I),
.I2(RIOB33_X105Y157_IOB_X1Y157_I),
.I3(CLBLL_L_X2Y134_SLICE_X0Y134_BO6),
.I4(LIOB33_X0Y151_IOB_X0Y152_I),
.I5(LIOB33_X0Y5_IOB_X0Y6_I),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_AO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_DO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_CO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_BO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_AO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_DO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_CO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_BO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555755555557)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_ALUT (
.I0(LIOB33_X0Y209_IOB_X0Y209_I),
.I1(LIOB33_X0Y161_IOB_X0Y162_I),
.I2(LIOB33_X0Y207_IOB_X0Y208_I),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I4(LIOB33_X0Y163_IOB_X0Y164_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_AO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_DO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_CO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_BO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_AO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he000e00000000000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_DLUT (
.I0(LIOB33_X0Y133_IOB_X0Y134_I),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I2(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I3(LIOB33_X0Y207_IOB_X0Y207_I),
.I4(1'b1),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_DO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f4f40000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_CLUT (
.I0(CLBLL_L_X2Y142_SLICE_X0Y142_AO6),
.I1(CLBLL_L_X2Y150_SLICE_X0Y150_AO6),
.I2(LIOB33_X0Y59_IOB_X0Y59_I),
.I3(1'b1),
.I4(CLBLL_L_X2Y142_SLICE_X0Y142_DO6),
.I5(CLBLL_L_X2Y142_SLICE_X0Y142_BO6),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_CO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_BLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(LIOB33_X0Y135_IOB_X0Y136_I),
.I3(LIOB33_X0Y119_IOB_X0Y119_I),
.I4(LIOB33_X0Y141_IOB_X0Y142_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_BO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffff)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_ALUT (
.I0(CLBLL_L_X2Y145_SLICE_X0Y145_DO6),
.I1(LIOB33_X0Y195_IOB_X0Y196_I),
.I2(LIOB33_X0Y139_IOB_X0Y140_I),
.I3(LIOB33_X0Y187_IOB_X0Y188_I),
.I4(CLBLL_L_X2Y131_SLICE_X0Y131_AO6),
.I5(LIOB33_X0Y89_IOB_X0Y89_I),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_AO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_DO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_CO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_BO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_AO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffefffe)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_DLUT (
.I0(LIOB33_X0Y145_IOB_X0Y145_I),
.I1(LIOB33_X0Y141_IOB_X0Y141_I),
.I2(LIOB33_X0Y181_IOB_X0Y181_I),
.I3(LIOB33_X0Y137_IOB_X0Y137_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_DO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc88cc8800000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I2(1'b1),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(1'b1),
.I5(LIOB33_X0Y205_IOB_X0Y206_I),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_CO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8f88888888888)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_BLUT (
.I0(LIOB33_X0Y139_IOB_X0Y140_I),
.I1(LIOB33_X0Y177_IOB_X0Y177_I),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(LIOB33_X0Y205_IOB_X0Y206_I),
.I4(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_BO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff80ff00)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_ALUT (
.I0(LIOB33_X0Y141_IOB_X0Y141_I),
.I1(LIOB33_X0Y141_IOB_X0Y142_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y145_SLICE_X0Y145_BO6),
.I4(LIOB33_X0Y145_IOB_X0Y145_I),
.I5(CLBLL_L_X2Y145_SLICE_X0Y145_CO6),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_AO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_DO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_CO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_BO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_AO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffff0000ffff)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y153_IOB_X0Y153_I),
.I3(1'b1),
.I4(LIOB33_X0Y129_IOB_X0Y130_I),
.I5(LIOB33_X0Y25_IOB_X0Y26_I),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccd00000005)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_ALUT (
.I0(LIOB33_X0Y155_IOB_X0Y156_I),
.I1(CLBLL_L_X2Y103_SLICE_X0Y103_BO6),
.I2(CLBLL_L_X2Y134_SLICE_X0Y134_CO6),
.I3(LIOB33_X0Y163_IOB_X0Y164_I),
.I4(LIOB33_X0Y161_IOB_X0Y162_I),
.I5(LIOB33_X0Y205_IOB_X0Y206_I),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff55550500)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_DLUT (
.I0(CLBLL_L_X2Y148_SLICE_X0Y148_AO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y149_SLICE_X0Y149_BO6),
.I3(CLBLL_L_X2Y149_SLICE_X0Y149_CO6),
.I4(CLBLL_L_X2Y149_SLICE_X0Y149_DO6),
.I5(CLBLL_L_X2Y148_SLICE_X0Y148_BO6),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000033300001333)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_CLUT (
.I0(LIOB33_X0Y139_IOB_X0Y139_I),
.I1(LIOB33_X0Y205_IOB_X0Y206_I),
.I2(CLBLL_L_X2Y103_SLICE_X1Y103_BO6),
.I3(LIOB33_X0Y181_IOB_X0Y182_I),
.I4(CLBLL_L_X2Y103_SLICE_X0Y103_BO6),
.I5(CLBLL_L_X2Y103_SLICE_X0Y103_AO6),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaa2a2a0)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_BLUT (
.I0(CLBLL_L_X2Y149_SLICE_X1Y149_AO5),
.I1(CLBLL_L_X2Y192_SLICE_X0Y192_DO6),
.I2(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I5(CLBLL_L_X2Y148_SLICE_X0Y148_CO6),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0cffffff5d)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_ALUT (
.I0(CLBLL_L_X2Y149_SLICE_X1Y149_AO5),
.I1(CLBLL_L_X2Y189_SLICE_X0Y189_CO6),
.I2(LIOB33_X0Y227_IOB_X0Y227_I),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I5(CLBLL_L_X2Y148_SLICE_X0Y148_CO6),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33a0a03333a0a0)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_DLUT (
.I0(CLBLL_L_X2Y193_SLICE_X0Y193_AO6),
.I1(CLBLL_L_X2Y149_SLICE_X1Y149_AO6),
.I2(CLBLL_L_X2Y149_SLICE_X1Y149_BO6),
.I3(1'b1),
.I4(LIOB33_X0Y227_IOB_X0Y227_I),
.I5(LIOB33_X0Y161_IOB_X0Y161_I),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_DO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefafce0affffcc00)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_CLUT (
.I0(CLBLL_L_X2Y149_SLICE_X0Y149_AO6),
.I1(CLBLL_L_X2Y149_SLICE_X1Y149_CO6),
.I2(CLBLL_L_X2Y150_SLICE_X0Y150_BO6),
.I3(CLBLL_L_X2Y210_SLICE_X0Y210_BO6),
.I4(CLBLL_L_X2Y208_SLICE_X0Y208_BO6),
.I5(CLBLL_L_X2Y149_SLICE_X1Y149_AO6),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_CO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003f0f33003b0a)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_BLUT (
.I0(LIOB33_X0Y141_IOB_X0Y141_I),
.I1(CLBLL_L_X2Y149_SLICE_X1Y149_BO6),
.I2(CLBLL_L_X2Y149_SLICE_X1Y149_AO6),
.I3(CLBLL_L_X2Y193_SLICE_X0Y193_DO6),
.I4(CLBLL_L_X2Y210_SLICE_X0Y210_BO6),
.I5(LIOB33_X0Y159_IOB_X0Y159_I),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_BO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0ffffffee)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_ALUT (
.I0(LIOB33_X0Y159_IOB_X0Y159_I),
.I1(LIOB33_X0Y157_IOB_X0Y157_I),
.I2(LIOB33_X0Y139_IOB_X0Y140_I),
.I3(LIOB33_X0Y161_IOB_X0Y161_I),
.I4(LIOB33_X0Y159_IOB_X0Y160_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_AO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_DO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddffdfdfdfff)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_CLUT (
.I0(LIOB33_X0Y181_IOB_X0Y182_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_BO6),
.I2(LIOB33_X0Y141_IOB_X0Y141_I),
.I3(CLBLL_L_X2Y103_SLICE_X0Y103_AO6),
.I4(LIOB33_X0Y139_IOB_X0Y139_I),
.I5(LIOB33_X0Y159_IOB_X0Y159_I),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_CO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcdffffcdffffff)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_BLUT (
.I0(LIOB33_X0Y141_IOB_X0Y142_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_BO6),
.I2(LIOB33_X0Y159_IOB_X0Y160_I),
.I3(CLBLL_L_X2Y103_SLICE_X0Y103_AO6),
.I4(LIOB33_X0Y181_IOB_X0Y182_I),
.I5(LIOB33_X0Y139_IOB_X0Y139_I),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_BO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddffff3377ffff)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_ALUT (
.I0(LIOB33_X0Y139_IOB_X0Y139_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_BO6),
.I2(1'b1),
.I3(CLBLL_L_X2Y103_SLICE_X0Y103_AO6),
.I4(LIOB33_X0Y181_IOB_X0Y182_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_AO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_DO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h02020202aaaaaaaa)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_CLUT (
.I0(LIOB33_X0Y133_IOB_X0Y133_I),
.I1(LIOB33_X0Y127_IOB_X0Y128_I),
.I2(CLBLL_L_X2Y193_SLICE_X0Y193_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y189_SLICE_X0Y189_BO6),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_CO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff8fffff88888888)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_BLUT (
.I0(LIOB33_X0Y155_IOB_X0Y156_I),
.I1(LIOB33_X0Y137_IOB_X0Y137_I),
.I2(LIOB33_X0Y135_IOB_X0Y136_I),
.I3(CLBLL_L_X2Y189_SLICE_X0Y189_BO6),
.I4(LIOB33_X0Y205_IOB_X0Y206_I),
.I5(CLBLL_L_X2Y193_SLICE_X0Y193_CO6),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_BO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee00eeee0e000e0e)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_ALUT (
.I0(CLBLL_L_X2Y193_SLICE_X0Y193_CO6),
.I1(LIOB33_X0Y137_IOB_X0Y137_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y189_SLICE_X0Y189_BO6),
.I4(LIOB33_X0Y135_IOB_X0Y136_I),
.I5(CLBLL_L_X2Y189_SLICE_X0Y189_CO6),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_AO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_DO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_CO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_BO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_AO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_DO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0f0f0a0a0f0f)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_CLUT (
.I0(CLBLL_L_X2Y151_SLICE_X0Y151_AO6),
.I1(1'b1),
.I2(LIOB33_X0Y179_IOB_X0Y180_I),
.I3(1'b1),
.I4(CLBLL_L_X2Y187_SLICE_X0Y187_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00400040f0f0f0f0)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_BLUT (
.I0(CLBLL_L_X2Y193_SLICE_X0Y193_CO6),
.I1(CLBLL_L_X2Y187_SLICE_X0Y187_BO6),
.I2(LIOB33_X0Y133_IOB_X0Y133_I),
.I3(LIOB33_X0Y127_IOB_X0Y128_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y210_SLICE_X0Y210_CO6),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_BO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff7)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_ALUT (
.I0(CLBLL_L_X2Y193_SLICE_X0Y193_CO6),
.I1(CLBLL_L_X2Y193_SLICE_X0Y193_AO6),
.I2(CLBLL_L_X2Y208_SLICE_X0Y208_BO6),
.I3(CLBLL_L_X2Y189_SLICE_X0Y189_BO6),
.I4(CLBLL_L_X2Y210_SLICE_X0Y210_BO6),
.I5(CLBLL_L_X2Y210_SLICE_X0Y210_CO6),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_AO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_DO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_CO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_BO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_AO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_DO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_CO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffff7f7fffff)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_BLUT (
.I0(LIOB33_X0Y207_IOB_X0Y208_I),
.I1(LIOB33_X0Y161_IOB_X0Y161_I),
.I2(LIOB33_X0Y209_IOB_X0Y209_I),
.I3(1'b1),
.I4(LIOB33_X0Y159_IOB_X0Y160_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_BO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0000000a00000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_ALUT (
.I0(LIOB33_X0Y155_IOB_X0Y156_I),
.I1(1'b1),
.I2(LIOB33_X0Y157_IOB_X0Y157_I),
.I3(CLBLL_L_X2Y154_SLICE_X0Y154_BO6),
.I4(LIOB33_X0Y159_IOB_X0Y159_I),
.I5(LIOB33_X0Y177_IOB_X0Y178_I),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_AO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_DO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_CO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y165_SLICE_X0Y165_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y165_SLICE_X0Y165_DO5),
.O6(CLBLL_L_X2Y165_SLICE_X0Y165_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c00000)
  ) CLBLL_L_X2Y165_SLICE_X0Y165_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y137_IOB_X0Y137_I),
.I2(LIOB33_X0Y135_IOB_X0Y136_I),
.I3(1'b1),
.I4(LIOB33_X0Y173_IOB_X0Y174_I),
.I5(LIOB33_X0Y175_IOB_X0Y175_I),
.O5(CLBLL_L_X2Y165_SLICE_X0Y165_CO5),
.O6(CLBLL_L_X2Y165_SLICE_X0Y165_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaa0a0aaaa)
  ) CLBLL_L_X2Y165_SLICE_X0Y165_BLUT (
.I0(LIOB33_X0Y15_IOB_X0Y15_I),
.I1(1'b1),
.I2(CLBLL_L_X2Y170_SLICE_X0Y170_AO6),
.I3(1'b1),
.I4(CLBLL_L_X2Y165_SLICE_X0Y165_AO6),
.I5(CLBLL_L_X2Y165_SLICE_X0Y165_CO6),
.O5(CLBLL_L_X2Y165_SLICE_X0Y165_BO5),
.O6(CLBLL_L_X2Y165_SLICE_X0Y165_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000057ff57ff57ff)
  ) CLBLL_L_X2Y165_SLICE_X0Y165_ALUT (
.I0(LIOB33_X0Y173_IOB_X0Y174_I),
.I1(LIOB33_X0Y135_IOB_X0Y136_I),
.I2(LIOB33_X0Y137_IOB_X0Y137_I),
.I3(LIOB33_X0Y175_IOB_X0Y175_I),
.I4(LIOB33_X0Y167_IOB_X0Y168_I),
.I5(LIOB33_X0Y165_IOB_X0Y166_I),
.O5(CLBLL_L_X2Y165_SLICE_X0Y165_AO5),
.O6(CLBLL_L_X2Y165_SLICE_X0Y165_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y165_SLICE_X1Y165_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y165_SLICE_X1Y165_DO5),
.O6(CLBLL_L_X2Y165_SLICE_X1Y165_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y165_SLICE_X1Y165_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y165_SLICE_X1Y165_CO5),
.O6(CLBLL_L_X2Y165_SLICE_X1Y165_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y165_SLICE_X1Y165_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y165_SLICE_X1Y165_BO5),
.O6(CLBLL_L_X2Y165_SLICE_X1Y165_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y165_SLICE_X1Y165_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y165_SLICE_X1Y165_AO5),
.O6(CLBLL_L_X2Y165_SLICE_X1Y165_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y170_SLICE_X0Y170_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y170_SLICE_X0Y170_DO5),
.O6(CLBLL_L_X2Y170_SLICE_X0Y170_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y170_SLICE_X0Y170_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y170_SLICE_X0Y170_CO5),
.O6(CLBLL_L_X2Y170_SLICE_X0Y170_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y170_SLICE_X0Y170_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y170_SLICE_X0Y170_BO5),
.O6(CLBLL_L_X2Y170_SLICE_X0Y170_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0000000a0000000)
  ) CLBLL_L_X2Y170_SLICE_X0Y170_ALUT (
.I0(LIOB33_X0Y171_IOB_X0Y172_I),
.I1(1'b1),
.I2(LIOB33_X0Y173_IOB_X0Y173_I),
.I3(LIOB33_X0Y169_IOB_X0Y169_I),
.I4(LIOB33_X0Y169_IOB_X0Y170_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y170_SLICE_X0Y170_AO5),
.O6(CLBLL_L_X2Y170_SLICE_X0Y170_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y170_SLICE_X1Y170_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y170_SLICE_X1Y170_DO5),
.O6(CLBLL_L_X2Y170_SLICE_X1Y170_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y170_SLICE_X1Y170_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y170_SLICE_X1Y170_CO5),
.O6(CLBLL_L_X2Y170_SLICE_X1Y170_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y170_SLICE_X1Y170_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y170_SLICE_X1Y170_BO5),
.O6(CLBLL_L_X2Y170_SLICE_X1Y170_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y170_SLICE_X1Y170_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y170_SLICE_X1Y170_AO5),
.O6(CLBLL_L_X2Y170_SLICE_X1Y170_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y187_SLICE_X0Y187_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y187_SLICE_X0Y187_DO5),
.O6(CLBLL_L_X2Y187_SLICE_X0Y187_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y187_SLICE_X0Y187_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y187_SLICE_X0Y187_CO5),
.O6(CLBLL_L_X2Y187_SLICE_X0Y187_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0e0c0f2e0)
  ) CLBLL_L_X2Y187_SLICE_X0Y187_BLUT (
.I0(CLBLL_L_X2Y189_SLICE_X0Y189_DO6),
.I1(LIOB33_X0Y153_IOB_X0Y154_I),
.I2(CLBLL_L_X2Y192_SLICE_X0Y192_AO6),
.I3(CLBLL_L_X2Y194_SLICE_X0Y194_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLL_L_X2Y187_SLICE_X0Y187_BO5),
.O6(CLBLL_L_X2Y187_SLICE_X0Y187_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000005500550055)
  ) CLBLL_L_X2Y187_SLICE_X0Y187_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y187_SLICE_X0Y187_AO5),
.O6(CLBLL_L_X2Y187_SLICE_X0Y187_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y187_SLICE_X1Y187_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y187_SLICE_X1Y187_DO5),
.O6(CLBLL_L_X2Y187_SLICE_X1Y187_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y187_SLICE_X1Y187_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y187_SLICE_X1Y187_CO5),
.O6(CLBLL_L_X2Y187_SLICE_X1Y187_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y187_SLICE_X1Y187_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y187_SLICE_X1Y187_BO5),
.O6(CLBLL_L_X2Y187_SLICE_X1Y187_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y187_SLICE_X1Y187_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y187_SLICE_X1Y187_AO5),
.O6(CLBLL_L_X2Y187_SLICE_X1Y187_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001010101)
  ) CLBLL_L_X2Y189_SLICE_X0Y189_DLUT (
.I0(LIOB33_X0Y233_IOB_X0Y234_I),
.I1(LIOB33_X0Y189_IOB_X0Y189_I),
.I2(LIOB33_X0Y221_IOB_X0Y222_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_SING_X0Y199_IOB_X0Y199_I),
.O5(CLBLL_L_X2Y189_SLICE_X0Y189_DO5),
.O6(CLBLL_L_X2Y189_SLICE_X0Y189_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000f000f000e)
  ) CLBLL_L_X2Y189_SLICE_X0Y189_CLUT (
.I0(LIOB33_X0Y233_IOB_X0Y234_I),
.I1(LIOB33_X0Y189_IOB_X0Y189_I),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(LIOB33_X0Y153_IOB_X0Y154_I),
.I4(LIOB33_X0Y221_IOB_X0Y222_I),
.I5(LIOB33_SING_X0Y199_IOB_X0Y199_I),
.O5(CLBLL_L_X2Y189_SLICE_X0Y189_CO5),
.O6(CLBLL_L_X2Y189_SLICE_X0Y189_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055555554)
  ) CLBLL_L_X2Y189_SLICE_X0Y189_BLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(LIOB33_X0Y229_IOB_X0Y229_I),
.I2(LIOB33_X0Y183_IOB_X0Y183_I),
.I3(LIOB33_X0Y193_IOB_X0Y194_I),
.I4(LIOB33_X0Y215_IOB_X0Y216_I),
.I5(LIOB33_X0Y153_IOB_X0Y154_I),
.O5(CLBLL_L_X2Y189_SLICE_X0Y189_BO5),
.O6(CLBLL_L_X2Y189_SLICE_X0Y189_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffd55555555)
  ) CLBLL_L_X2Y189_SLICE_X0Y189_ALUT (
.I0(LIOB33_X0Y131_IOB_X0Y132_I),
.I1(LIOB33_X0Y229_IOB_X0Y229_I),
.I2(LIOB33_X0Y183_IOB_X0Y183_I),
.I3(LIOB33_X0Y193_IOB_X0Y194_I),
.I4(LIOB33_X0Y215_IOB_X0Y216_I),
.I5(CLBLL_L_X2Y187_SLICE_X0Y187_AO5),
.O5(CLBLL_L_X2Y189_SLICE_X0Y189_AO5),
.O6(CLBLL_L_X2Y189_SLICE_X0Y189_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y189_SLICE_X1Y189_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y189_SLICE_X1Y189_DO5),
.O6(CLBLL_L_X2Y189_SLICE_X1Y189_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y189_SLICE_X1Y189_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y189_SLICE_X1Y189_CO5),
.O6(CLBLL_L_X2Y189_SLICE_X1Y189_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y189_SLICE_X1Y189_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y189_SLICE_X1Y189_BO5),
.O6(CLBLL_L_X2Y189_SLICE_X1Y189_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaaaaaab)
  ) CLBLL_L_X2Y189_SLICE_X1Y189_ALUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(LIOB33_SING_X0Y199_IOB_X0Y199_I),
.I2(LIOB33_X0Y189_IOB_X0Y189_I),
.I3(LIOB33_X0Y221_IOB_X0Y222_I),
.I4(LIOB33_X0Y233_IOB_X0Y234_I),
.I5(LIOB33_X0Y153_IOB_X0Y154_I),
.O5(CLBLL_L_X2Y189_SLICE_X1Y189_AO5),
.O6(CLBLL_L_X2Y189_SLICE_X1Y189_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00ff01ff)
  ) CLBLL_L_X2Y192_SLICE_X0Y192_DLUT (
.I0(LIOB33_X0Y231_IOB_X0Y231_I),
.I1(LIOB33_X0Y185_IOB_X0Y185_I),
.I2(LIOB33_X0Y197_IOB_X0Y197_I),
.I3(CLBLL_L_X2Y187_SLICE_X0Y187_AO5),
.I4(LIOB33_X0Y219_IOB_X0Y219_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X2Y192_SLICE_X0Y192_DO5),
.O6(CLBLL_L_X2Y192_SLICE_X0Y192_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003300330032)
  ) CLBLL_L_X2Y192_SLICE_X0Y192_CLUT (
.I0(LIOB33_X0Y191_IOB_X0Y192_I),
.I1(LIOB33_X0Y153_IOB_X0Y154_I),
.I2(LIOB33_X0Y213_IOB_X0Y214_I),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(LIOB33_X0Y237_IOB_X0Y238_I),
.I5(LIOB33_X0Y225_IOB_X0Y226_I),
.O5(CLBLL_L_X2Y192_SLICE_X0Y192_CO5),
.O6(CLBLL_L_X2Y192_SLICE_X0Y192_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000002aaaaaaaa)
  ) CLBLL_L_X2Y192_SLICE_X0Y192_BLUT (
.I0(LIOB33_X0Y133_IOB_X0Y133_I),
.I1(LIOB33_X0Y237_IOB_X0Y238_I),
.I2(LIOB33_X0Y191_IOB_X0Y192_I),
.I3(LIOB33_X0Y225_IOB_X0Y226_I),
.I4(LIOB33_X0Y213_IOB_X0Y214_I),
.I5(CLBLL_L_X2Y210_SLICE_X0Y210_BO6),
.O5(CLBLL_L_X2Y192_SLICE_X0Y192_BO5),
.O6(CLBLL_L_X2Y192_SLICE_X0Y192_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00ff01)
  ) CLBLL_L_X2Y192_SLICE_X0Y192_ALUT (
.I0(LIOB33_X0Y219_IOB_X0Y219_I),
.I1(LIOB33_X0Y231_IOB_X0Y231_I),
.I2(LIOB33_X0Y185_IOB_X0Y185_I),
.I3(LIOB33_X0Y153_IOB_X0Y154_I),
.I4(LIOB33_X0Y197_IOB_X0Y197_I),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLL_L_X2Y192_SLICE_X0Y192_AO5),
.O6(CLBLL_L_X2Y192_SLICE_X0Y192_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y192_SLICE_X1Y192_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y192_SLICE_X1Y192_DO5),
.O6(CLBLL_L_X2Y192_SLICE_X1Y192_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y192_SLICE_X1Y192_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y192_SLICE_X1Y192_CO5),
.O6(CLBLL_L_X2Y192_SLICE_X1Y192_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y192_SLICE_X1Y192_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y192_SLICE_X1Y192_BO5),
.O6(CLBLL_L_X2Y192_SLICE_X1Y192_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y192_SLICE_X1Y192_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y192_SLICE_X1Y192_AO5),
.O6(CLBLL_L_X2Y192_SLICE_X1Y192_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300330033003200)
  ) CLBLL_L_X2Y193_SLICE_X0Y193_DLUT (
.I0(LIOB33_X0Y189_IOB_X0Y190_I),
.I1(LIOB33_X0Y227_IOB_X0Y227_I),
.I2(LIOB33_X0Y223_IOB_X0Y223_I),
.I3(CLBLL_L_X2Y187_SLICE_X0Y187_AO5),
.I4(LIOB33_X0Y211_IOB_X0Y211_I),
.I5(LIOB33_X0Y235_IOB_X0Y235_I),
.O5(CLBLL_L_X2Y193_SLICE_X0Y193_DO5),
.O6(CLBLL_L_X2Y193_SLICE_X0Y193_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccffccffcd)
  ) CLBLL_L_X2Y193_SLICE_X0Y193_CLUT (
.I0(LIOB33_X0Y191_IOB_X0Y192_I),
.I1(LIOB33_X0Y153_IOB_X0Y154_I),
.I2(LIOB33_X0Y213_IOB_X0Y214_I),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(LIOB33_X0Y237_IOB_X0Y238_I),
.I5(LIOB33_X0Y225_IOB_X0Y226_I),
.O5(CLBLL_L_X2Y193_SLICE_X0Y193_CO5),
.O6(CLBLL_L_X2Y193_SLICE_X0Y193_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h222222222222222a)
  ) CLBLL_L_X2Y193_SLICE_X0Y193_BLUT (
.I0(LIOB33_X0Y133_IOB_X0Y133_I),
.I1(CLBLL_L_X2Y208_SLICE_X0Y208_BO6),
.I2(LIOB33_X0Y211_IOB_X0Y211_I),
.I3(LIOB33_X0Y223_IOB_X0Y223_I),
.I4(LIOB33_X0Y189_IOB_X0Y190_I),
.I5(LIOB33_X0Y235_IOB_X0Y235_I),
.O5(CLBLL_L_X2Y193_SLICE_X0Y193_BO5),
.O6(CLBLL_L_X2Y193_SLICE_X0Y193_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaaffffaaab)
  ) CLBLL_L_X2Y193_SLICE_X0Y193_ALUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(LIOB33_X0Y211_IOB_X0Y211_I),
.I2(LIOB33_X0Y189_IOB_X0Y190_I),
.I3(LIOB33_X0Y223_IOB_X0Y223_I),
.I4(LIOB33_X0Y153_IOB_X0Y154_I),
.I5(LIOB33_X0Y235_IOB_X0Y235_I),
.O5(CLBLL_L_X2Y193_SLICE_X0Y193_AO5),
.O6(CLBLL_L_X2Y193_SLICE_X0Y193_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y193_SLICE_X1Y193_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y193_SLICE_X1Y193_DO5),
.O6(CLBLL_L_X2Y193_SLICE_X1Y193_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y193_SLICE_X1Y193_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y193_SLICE_X1Y193_CO5),
.O6(CLBLL_L_X2Y193_SLICE_X1Y193_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y193_SLICE_X1Y193_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y193_SLICE_X1Y193_BO5),
.O6(CLBLL_L_X2Y193_SLICE_X1Y193_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y193_SLICE_X1Y193_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y193_SLICE_X1Y193_AO5),
.O6(CLBLL_L_X2Y193_SLICE_X1Y193_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y194_SLICE_X0Y194_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y194_SLICE_X0Y194_DO5),
.O6(CLBLL_L_X2Y194_SLICE_X0Y194_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y194_SLICE_X0Y194_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y194_SLICE_X0Y194_CO5),
.O6(CLBLL_L_X2Y194_SLICE_X0Y194_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000303)
  ) CLBLL_L_X2Y194_SLICE_X0Y194_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y219_IOB_X0Y220_I),
.I2(LIOB33_X0Y185_IOB_X0Y186_I),
.I3(1'b1),
.I4(LIOB33_X0Y231_IOB_X0Y232_I),
.I5(LIOB33_X0Y197_IOB_X0Y198_I),
.O5(CLBLL_L_X2Y194_SLICE_X0Y194_BO5),
.O6(CLBLL_L_X2Y194_SLICE_X0Y194_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaaaaaab)
  ) CLBLL_L_X2Y194_SLICE_X0Y194_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(LIOB33_X0Y219_IOB_X0Y220_I),
.I2(LIOB33_X0Y185_IOB_X0Y186_I),
.I3(LIOB33_X0Y197_IOB_X0Y198_I),
.I4(LIOB33_X0Y231_IOB_X0Y232_I),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLL_L_X2Y194_SLICE_X0Y194_AO5),
.O6(CLBLL_L_X2Y194_SLICE_X0Y194_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y194_SLICE_X1Y194_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y194_SLICE_X1Y194_DO5),
.O6(CLBLL_L_X2Y194_SLICE_X1Y194_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y194_SLICE_X1Y194_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y194_SLICE_X1Y194_CO5),
.O6(CLBLL_L_X2Y194_SLICE_X1Y194_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y194_SLICE_X1Y194_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y194_SLICE_X1Y194_BO5),
.O6(CLBLL_L_X2Y194_SLICE_X1Y194_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y194_SLICE_X1Y194_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y194_SLICE_X1Y194_AO5),
.O6(CLBLL_L_X2Y194_SLICE_X1Y194_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y208_SLICE_X0Y208_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y208_SLICE_X0Y208_DO5),
.O6(CLBLL_L_X2Y208_SLICE_X0Y208_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y208_SLICE_X0Y208_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y208_SLICE_X0Y208_CO5),
.O6(CLBLL_L_X2Y208_SLICE_X0Y208_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033333332)
  ) CLBLL_L_X2Y208_SLICE_X0Y208_BLUT (
.I0(LIOB33_X0Y213_IOB_X0Y213_I),
.I1(LIOB33_X0Y153_IOB_X0Y154_I),
.I2(LIOB33_X0Y191_IOB_X0Y191_I),
.I3(LIOB33_X0Y237_IOB_X0Y237_I),
.I4(LIOB33_X0Y225_IOB_X0Y225_I),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLL_L_X2Y208_SLICE_X0Y208_BO5),
.O6(CLBLL_L_X2Y208_SLICE_X0Y208_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcccccccd)
  ) CLBLL_L_X2Y208_SLICE_X0Y208_ALUT (
.I0(LIOB33_X0Y213_IOB_X0Y213_I),
.I1(LIOB33_X0Y153_IOB_X0Y154_I),
.I2(LIOB33_X0Y225_IOB_X0Y225_I),
.I3(LIOB33_X0Y237_IOB_X0Y237_I),
.I4(LIOB33_X0Y191_IOB_X0Y191_I),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLL_L_X2Y208_SLICE_X0Y208_AO5),
.O6(CLBLL_L_X2Y208_SLICE_X0Y208_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y208_SLICE_X1Y208_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y208_SLICE_X1Y208_DO5),
.O6(CLBLL_L_X2Y208_SLICE_X1Y208_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y208_SLICE_X1Y208_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y208_SLICE_X1Y208_CO5),
.O6(CLBLL_L_X2Y208_SLICE_X1Y208_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y208_SLICE_X1Y208_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y208_SLICE_X1Y208_BO5),
.O6(CLBLL_L_X2Y208_SLICE_X1Y208_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y208_SLICE_X1Y208_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y208_SLICE_X1Y208_AO5),
.O6(CLBLL_L_X2Y208_SLICE_X1Y208_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y210_SLICE_X0Y210_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y210_SLICE_X0Y210_DO5),
.O6(CLBLL_L_X2Y210_SLICE_X0Y210_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003300330032)
  ) CLBLL_L_X2Y210_SLICE_X0Y210_CLUT (
.I0(LIOB33_X0Y215_IOB_X0Y215_I),
.I1(LIOB33_X0Y153_IOB_X0Y154_I),
.I2(LIOB33_X0Y239_IOB_X0Y239_I),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(LIOB33_X0Y193_IOB_X0Y193_I),
.I5(LIOB33_X0Y227_IOB_X0Y228_I),
.O5(CLBLL_L_X2Y210_SLICE_X0Y210_CO5),
.O6(CLBLL_L_X2Y210_SLICE_X0Y210_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033333332)
  ) CLBLL_L_X2Y210_SLICE_X0Y210_BLUT (
.I0(LIOB33_X0Y211_IOB_X0Y212_I),
.I1(LIOB33_X0Y153_IOB_X0Y154_I),
.I2(LIOB33_X0Y209_IOB_X0Y210_I),
.I3(LIOB33_X0Y235_IOB_X0Y236_I),
.I4(LIOB33_X0Y223_IOB_X0Y224_I),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLL_L_X2Y210_SLICE_X0Y210_BO5),
.O6(CLBLL_L_X2Y210_SLICE_X0Y210_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00ff01)
  ) CLBLL_L_X2Y210_SLICE_X0Y210_ALUT (
.I0(LIOB33_X0Y211_IOB_X0Y212_I),
.I1(LIOB33_X0Y223_IOB_X0Y224_I),
.I2(LIOB33_X0Y209_IOB_X0Y210_I),
.I3(LIOB33_X0Y153_IOB_X0Y154_I),
.I4(LIOB33_X0Y235_IOB_X0Y236_I),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLL_L_X2Y210_SLICE_X0Y210_AO5),
.O6(CLBLL_L_X2Y210_SLICE_X0Y210_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y210_SLICE_X1Y210_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y210_SLICE_X1Y210_DO5),
.O6(CLBLL_L_X2Y210_SLICE_X1Y210_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y210_SLICE_X1Y210_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y210_SLICE_X1Y210_CO5),
.O6(CLBLL_L_X2Y210_SLICE_X1Y210_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y210_SLICE_X1Y210_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y210_SLICE_X1Y210_BO5),
.O6(CLBLL_L_X2Y210_SLICE_X1Y210_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y210_SLICE_X1Y210_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y210_SLICE_X1Y210_AO5),
.O6(CLBLL_L_X2Y210_SLICE_X1Y210_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y152_SLICE_X66Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y152_SLICE_X66Y152_DO5),
.O6(CLBLM_L_X44Y152_SLICE_X66Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y152_SLICE_X66Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y152_SLICE_X66Y152_CO5),
.O6(CLBLM_L_X44Y152_SLICE_X66Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y152_SLICE_X66Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y152_SLICE_X66Y152_BO5),
.O6(CLBLM_L_X44Y152_SLICE_X66Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefffaff55555555)
  ) CLBLM_L_X44Y152_SLICE_X66Y152_ALUT (
.I0(CLBLM_R_X47Y158_SLICE_X72Y158_BO6),
.I1(LIOB33_X0Y157_IOB_X0Y158_I),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(LIOB33_X0Y129_IOB_X0Y130_I),
.I4(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I5(1'b1),
.O5(CLBLM_L_X44Y152_SLICE_X66Y152_AO5),
.O6(CLBLM_L_X44Y152_SLICE_X66Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y152_SLICE_X67Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y152_SLICE_X67Y152_DO5),
.O6(CLBLM_L_X44Y152_SLICE_X67Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y152_SLICE_X67Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y152_SLICE_X67Y152_CO5),
.O6(CLBLM_L_X44Y152_SLICE_X67Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y152_SLICE_X67Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y152_SLICE_X67Y152_BO5),
.O6(CLBLM_L_X44Y152_SLICE_X67Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y152_SLICE_X67Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y152_SLICE_X67Y152_AO5),
.O6(CLBLM_L_X44Y152_SLICE_X67Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y158_SLICE_X66Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y158_SLICE_X66Y158_DO5),
.O6(CLBLM_L_X44Y158_SLICE_X66Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y158_SLICE_X66Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y158_SLICE_X66Y158_CO5),
.O6(CLBLM_L_X44Y158_SLICE_X66Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffff5f5f5f5f)
  ) CLBLM_L_X44Y158_SLICE_X66Y158_BLUT (
.I0(LIOB33_X0Y129_IOB_X0Y130_I),
.I1(LIOB33_X0Y125_IOB_X0Y125_I),
.I2(LIOB33_X0Y217_IOB_X0Y218_I),
.I3(CLBLM_R_X47Y158_SLICE_X72Y158_BO6),
.I4(LIOB33_X0Y179_IOB_X0Y179_I),
.I5(1'b1),
.O5(CLBLM_L_X44Y158_SLICE_X66Y158_BO5),
.O6(CLBLM_L_X44Y158_SLICE_X66Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0ffa0ffa0a0ffff)
  ) CLBLM_L_X44Y158_SLICE_X66Y158_ALUT (
.I0(LIOB33_X0Y129_IOB_X0Y130_I),
.I1(1'b1),
.I2(LIOB33_X0Y217_IOB_X0Y218_I),
.I3(LIOB33_X0Y165_IOB_X0Y165_I),
.I4(LIOB33_X0Y129_IOB_X0Y129_I),
.I5(1'b1),
.O5(CLBLM_L_X44Y158_SLICE_X66Y158_AO5),
.O6(CLBLM_L_X44Y158_SLICE_X66Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y158_SLICE_X67Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y158_SLICE_X67Y158_DO5),
.O6(CLBLM_L_X44Y158_SLICE_X67Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y158_SLICE_X67Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y158_SLICE_X67Y158_CO5),
.O6(CLBLM_L_X44Y158_SLICE_X67Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y158_SLICE_X67Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y158_SLICE_X67Y158_BO5),
.O6(CLBLM_L_X44Y158_SLICE_X67Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y158_SLICE_X67Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y158_SLICE_X67Y158_AO5),
.O6(CLBLM_L_X44Y158_SLICE_X67Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y145_SLICE_X72Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y145_SLICE_X72Y145_DO5),
.O6(CLBLM_R_X47Y145_SLICE_X72Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y145_SLICE_X72Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y145_SLICE_X72Y145_CO5),
.O6(CLBLM_R_X47Y145_SLICE_X72Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y145_SLICE_X72Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y145_SLICE_X72Y145_BO5),
.O6(CLBLM_R_X47Y145_SLICE_X72Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001010101)
  ) CLBLM_R_X47Y145_SLICE_X72Y145_ALUT (
.I0(LIOB33_X0Y217_IOB_X0Y217_I),
.I1(LIOB33_X0Y1_IOB_X0Y1_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y195_IOB_X0Y195_I),
.O5(CLBLM_R_X47Y145_SLICE_X72Y145_AO5),
.O6(CLBLM_R_X47Y145_SLICE_X72Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y145_SLICE_X73Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y145_SLICE_X73Y145_DO5),
.O6(CLBLM_R_X47Y145_SLICE_X73Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y145_SLICE_X73Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y145_SLICE_X73Y145_CO5),
.O6(CLBLM_R_X47Y145_SLICE_X73Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y145_SLICE_X73Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y145_SLICE_X73Y145_BO5),
.O6(CLBLM_R_X47Y145_SLICE_X73Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y145_SLICE_X73Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y145_SLICE_X73Y145_AO5),
.O6(CLBLM_R_X47Y145_SLICE_X73Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y158_SLICE_X72Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y158_SLICE_X72Y158_DO5),
.O6(CLBLM_R_X47Y158_SLICE_X72Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y158_SLICE_X72Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y158_SLICE_X72Y158_CO5),
.O6(CLBLM_R_X47Y158_SLICE_X72Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff0000f0fff0ff)
  ) CLBLM_R_X47Y158_SLICE_X72Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X47Y145_SLICE_X72Y145_AO6),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(CLBLM_R_X47Y158_SLICE_X72Y158_AO6),
.I5(LIOB33_X0Y165_IOB_X0Y165_I),
.O5(CLBLM_R_X47Y158_SLICE_X72Y158_BO5),
.O6(CLBLM_R_X47Y158_SLICE_X72Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000010)
  ) CLBLM_R_X47Y158_SLICE_X72Y158_ALUT (
.I0(LIOB33_X0Y229_IOB_X0Y230_I),
.I1(LIOB33_X0Y241_IOB_X0Y242_I),
.I2(CLBLM_R_X47Y145_SLICE_X72Y145_AO6),
.I3(LIOB33_X0Y183_IOB_X0Y184_I),
.I4(LIOB33_X0Y9_IOB_X0Y10_I),
.I5(1'b1),
.O5(CLBLM_R_X47Y158_SLICE_X72Y158_AO5),
.O6(CLBLM_R_X47Y158_SLICE_X72Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y158_SLICE_X73Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y158_SLICE_X73Y158_DO5),
.O6(CLBLM_R_X47Y158_SLICE_X73Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y158_SLICE_X73Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y158_SLICE_X73Y158_CO5),
.O6(CLBLM_R_X47Y158_SLICE_X73Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y158_SLICE_X73Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y158_SLICE_X73Y158_BO5),
.O6(CLBLM_R_X47Y158_SLICE_X73Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X47Y158_SLICE_X73Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X47Y158_SLICE_X73Y158_AO5),
.O6(CLBLM_R_X47Y158_SLICE_X73Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y133_SLICE_X88Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y133_SLICE_X88Y133_DO5),
.O6(CLBLM_R_X59Y133_SLICE_X88Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y133_SLICE_X88Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y133_SLICE_X88Y133_CO5),
.O6(CLBLM_R_X59Y133_SLICE_X88Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y133_SLICE_X88Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y133_SLICE_X88Y133_BO5),
.O6(CLBLM_R_X59Y133_SLICE_X88Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X59Y133_SLICE_X88Y133_ALUT (
.I0(CLBLL_L_X2Y134_SLICE_X0Y134_AO6),
.I1(CLBLM_R_X47Y158_SLICE_X72Y158_BO6),
.I2(CLBLL_L_X2Y165_SLICE_X0Y165_BO6),
.I3(CLBLL_L_X2Y145_SLICE_X0Y145_AO6),
.I4(CLBLL_L_X2Y154_SLICE_X0Y154_AO6),
.I5(CLBLL_L_X2Y151_SLICE_X0Y151_CO6),
.O5(CLBLM_R_X59Y133_SLICE_X88Y133_AO5),
.O6(CLBLM_R_X59Y133_SLICE_X88Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y133_SLICE_X89Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y133_SLICE_X89Y133_DO5),
.O6(CLBLM_R_X59Y133_SLICE_X89Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y133_SLICE_X89Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y133_SLICE_X89Y133_CO5),
.O6(CLBLM_R_X59Y133_SLICE_X89Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y133_SLICE_X89Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y133_SLICE_X89Y133_BO5),
.O6(CLBLM_R_X59Y133_SLICE_X89Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y133_SLICE_X89Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y133_SLICE_X89Y133_AO5),
.O6(CLBLM_R_X59Y133_SLICE_X89Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y159_SLICE_X88Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y159_SLICE_X88Y159_DO5),
.O6(CLBLM_R_X59Y159_SLICE_X88Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y159_SLICE_X88Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y159_SLICE_X88Y159_CO5),
.O6(CLBLM_R_X59Y159_SLICE_X88Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y159_SLICE_X88Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y159_SLICE_X88Y159_BO5),
.O6(CLBLM_R_X59Y159_SLICE_X88Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f5f5f5f5f)
  ) CLBLM_R_X59Y159_SLICE_X88Y159_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(1'b1),
.I2(LIOB33_X0Y239_IOB_X0Y240_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y159_SLICE_X88Y159_AO5),
.O6(CLBLM_R_X59Y159_SLICE_X88Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y159_SLICE_X89Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y159_SLICE_X89Y159_DO5),
.O6(CLBLM_R_X59Y159_SLICE_X89Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y159_SLICE_X89Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y159_SLICE_X89Y159_CO5),
.O6(CLBLM_R_X59Y159_SLICE_X89Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y159_SLICE_X89Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y159_SLICE_X89Y159_BO5),
.O6(CLBLM_R_X59Y159_SLICE_X89Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y159_SLICE_X89Y159_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y159_SLICE_X89Y159_AO5),
.O6(CLBLM_R_X59Y159_SLICE_X89Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y130_SLICE_X100Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y130_SLICE_X100Y130_DO5),
.O6(CLBLM_R_X67Y130_SLICE_X100Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y130_SLICE_X100Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y130_SLICE_X100Y130_CO5),
.O6(CLBLM_R_X67Y130_SLICE_X100Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y130_SLICE_X100Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y130_SLICE_X100Y130_BO5),
.O6(CLBLM_R_X67Y130_SLICE_X100Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X67Y130_SLICE_X100Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y165_SLICE_X0Y165_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y130_SLICE_X100Y130_AO5),
.O6(CLBLM_R_X67Y130_SLICE_X100Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y130_SLICE_X101Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y130_SLICE_X101Y130_DO5),
.O6(CLBLM_R_X67Y130_SLICE_X101Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y130_SLICE_X101Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y130_SLICE_X101Y130_CO5),
.O6(CLBLM_R_X67Y130_SLICE_X101Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y130_SLICE_X101Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y130_SLICE_X101Y130_BO5),
.O6(CLBLM_R_X67Y130_SLICE_X101Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X67Y130_SLICE_X101Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X67Y130_SLICE_X101Y130_AO5),
.O6(CLBLM_R_X67Y130_SLICE_X101Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y1_IOB_X0Y1_IBUF (
.I(LIOB33_X0Y1_IOB_X0Y1_IPAD),
.O(LIOB33_X0Y1_IOB_X0Y1_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y1_IOB_X0Y2_IBUF (
.I(LIOB33_X0Y1_IOB_X0Y2_IPAD),
.O(LIOB33_X0Y1_IOB_X0Y2_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y3_IOB_X0Y3_IBUF (
.I(LIOB33_X0Y3_IOB_X0Y3_IPAD),
.O(LIOB33_X0Y3_IOB_X0Y3_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y3_IOB_X0Y4_IBUF (
.I(LIOB33_X0Y3_IOB_X0Y4_IPAD),
.O(LIOB33_X0Y3_IOB_X0Y4_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y5_IOB_X0Y5_IBUF (
.I(LIOB33_X0Y5_IOB_X0Y5_IPAD),
.O(LIOB33_X0Y5_IOB_X0Y5_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y5_IOB_X0Y6_IBUF (
.I(LIOB33_X0Y5_IOB_X0Y6_IPAD),
.O(LIOB33_X0Y5_IOB_X0Y6_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y7_IOB_X0Y7_IBUF (
.I(LIOB33_X0Y7_IOB_X0Y7_IPAD),
.O(LIOB33_X0Y7_IOB_X0Y7_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y7_IOB_X0Y8_IBUF (
.I(LIOB33_X0Y7_IOB_X0Y8_IPAD),
.O(LIOB33_X0Y7_IOB_X0Y8_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y9_IOB_X0Y9_IBUF (
.I(LIOB33_X0Y9_IOB_X0Y9_IPAD),
.O(LIOB33_X0Y9_IOB_X0Y9_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y9_IOB_X0Y10_IBUF (
.I(LIOB33_X0Y9_IOB_X0Y10_IPAD),
.O(LIOB33_X0Y9_IOB_X0Y10_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(LIOB33_X0Y11_IOB_X0Y11_IPAD),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y11_IOB_X0Y12_IBUF (
.I(LIOB33_X0Y11_IOB_X0Y12_IPAD),
.O(LIOB33_X0Y11_IOB_X0Y12_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y13_IOB_X0Y13_IBUF (
.I(LIOB33_X0Y13_IOB_X0Y13_IPAD),
.O(LIOB33_X0Y13_IOB_X0Y13_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y13_IOB_X0Y14_IBUF (
.I(LIOB33_X0Y13_IOB_X0Y14_IPAD),
.O(LIOB33_X0Y13_IOB_X0Y14_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y15_IOB_X0Y15_IBUF (
.I(LIOB33_X0Y15_IOB_X0Y15_IPAD),
.O(LIOB33_X0Y15_IOB_X0Y15_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y15_IOB_X0Y16_IBUF (
.I(LIOB33_X0Y15_IOB_X0Y16_IPAD),
.O(LIOB33_X0Y15_IOB_X0Y16_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y17_IOB_X0Y17_IBUF (
.I(LIOB33_X0Y17_IOB_X0Y17_IPAD),
.O(LIOB33_X0Y17_IOB_X0Y17_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y17_IOB_X0Y18_IBUF (
.I(LIOB33_X0Y17_IOB_X0Y18_IPAD),
.O(LIOB33_X0Y17_IOB_X0Y18_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y19_IOB_X0Y19_IBUF (
.I(LIOB33_X0Y19_IOB_X0Y19_IPAD),
.O(LIOB33_X0Y19_IOB_X0Y19_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y19_IOB_X0Y20_IBUF (
.I(LIOB33_X0Y19_IOB_X0Y20_IPAD),
.O(LIOB33_X0Y19_IOB_X0Y20_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y21_IOB_X0Y21_IBUF (
.I(LIOB33_X0Y21_IOB_X0Y21_IPAD),
.O(LIOB33_X0Y21_IOB_X0Y21_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y21_IOB_X0Y22_IBUF (
.I(LIOB33_X0Y21_IOB_X0Y22_IPAD),
.O(LIOB33_X0Y21_IOB_X0Y22_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y23_IOB_X0Y23_IBUF (
.I(LIOB33_X0Y23_IOB_X0Y23_IPAD),
.O(LIOB33_X0Y23_IOB_X0Y23_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y23_IOB_X0Y24_IBUF (
.I(LIOB33_X0Y23_IOB_X0Y24_IPAD),
.O(LIOB33_X0Y23_IOB_X0Y24_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y25_IOB_X0Y25_IBUF (
.I(LIOB33_X0Y25_IOB_X0Y25_IPAD),
.O(LIOB33_X0Y25_IOB_X0Y25_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y25_IOB_X0Y26_IBUF (
.I(LIOB33_X0Y25_IOB_X0Y26_IPAD),
.O(LIOB33_X0Y25_IOB_X0Y26_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y27_IOB_X0Y27_IBUF (
.I(LIOB33_X0Y27_IOB_X0Y27_IPAD),
.O(LIOB33_X0Y27_IOB_X0Y27_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y27_IOB_X0Y28_IBUF (
.I(LIOB33_X0Y27_IOB_X0Y28_IPAD),
.O(LIOB33_X0Y27_IOB_X0Y28_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y80_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y80_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y81_IOB_X0Y81_IBUF (
.I(LIOB33_X0Y81_IOB_X0Y81_IPAD),
.O(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y81_IOB_X0Y82_IBUF (
.I(LIOB33_X0Y81_IOB_X0Y82_IPAD),
.O(LIOB33_X0Y81_IOB_X0Y82_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y83_IOB_X0Y83_IBUF (
.I(LIOB33_X0Y83_IOB_X0Y83_IPAD),
.O(LIOB33_X0Y83_IOB_X0Y83_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y83_IOB_X0Y84_IBUF (
.I(LIOB33_X0Y83_IOB_X0Y84_IPAD),
.O(LIOB33_X0Y83_IOB_X0Y84_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y85_IOB_X0Y85_IBUF (
.I(LIOB33_X0Y85_IOB_X0Y85_IPAD),
.O(LIOB33_X0Y85_IOB_X0Y85_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y85_IOB_X0Y86_IBUF (
.I(LIOB33_X0Y85_IOB_X0Y86_IPAD),
.O(LIOB33_X0Y85_IOB_X0Y86_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y87_IOB_X0Y87_IBUF (
.I(LIOB33_X0Y87_IOB_X0Y87_IPAD),
.O(LIOB33_X0Y87_IOB_X0Y87_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y87_IOB_X0Y88_IBUF (
.I(LIOB33_X0Y87_IOB_X0Y88_IPAD),
.O(LIOB33_X0Y87_IOB_X0Y88_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y89_IOB_X0Y89_IBUF (
.I(LIOB33_X0Y89_IOB_X0Y89_IPAD),
.O(LIOB33_X0Y89_IOB_X0Y89_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y89_IOB_X0Y90_IBUF (
.I(LIOB33_X0Y89_IOB_X0Y90_IPAD),
.O(LIOB33_X0Y89_IOB_X0Y90_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y91_IOB_X0Y91_IBUF (
.I(LIOB33_X0Y91_IOB_X0Y91_IPAD),
.O(LIOB33_X0Y91_IOB_X0Y91_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y91_IOB_X0Y92_IBUF (
.I(LIOB33_X0Y91_IOB_X0Y92_IPAD),
.O(LIOB33_X0Y91_IOB_X0Y92_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y93_IOB_X0Y93_IBUF (
.I(LIOB33_X0Y93_IOB_X0Y93_IPAD),
.O(LIOB33_X0Y93_IOB_X0Y93_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y93_IOB_X0Y94_IBUF (
.I(LIOB33_X0Y93_IOB_X0Y94_IPAD),
.O(LIOB33_X0Y93_IOB_X0Y94_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y95_IOB_X0Y95_IBUF (
.I(LIOB33_X0Y95_IOB_X0Y95_IPAD),
.O(LIOB33_X0Y95_IOB_X0Y95_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y95_IOB_X0Y96_IBUF (
.I(LIOB33_X0Y95_IOB_X0Y96_IPAD),
.O(LIOB33_X0Y95_IOB_X0Y96_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y97_IOB_X0Y97_IBUF (
.I(LIOB33_X0Y97_IOB_X0Y97_IPAD),
.O(LIOB33_X0Y97_IOB_X0Y97_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y97_IOB_X0Y98_IBUF (
.I(LIOB33_X0Y97_IOB_X0Y98_IPAD),
.O(LIOB33_X0Y97_IOB_X0Y98_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y119_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y119_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y120_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y120_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y121_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y121_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y122_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y124_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y125_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y126_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y127_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y128_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y129_IOB_X0Y129_IBUF (
.I(LIOB33_X0Y129_IOB_X0Y129_IPAD),
.O(LIOB33_X0Y129_IOB_X0Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y129_IOB_X0Y130_IBUF (
.I(LIOB33_X0Y129_IOB_X0Y130_IPAD),
.O(LIOB33_X0Y129_IOB_X0Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y131_IOB_X0Y131_IBUF (
.I(LIOB33_X0Y131_IOB_X0Y131_IPAD),
.O(LIOB33_X0Y131_IOB_X0Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y131_IOB_X0Y132_IBUF (
.I(LIOB33_X0Y131_IOB_X0Y132_IPAD),
.O(LIOB33_X0Y131_IOB_X0Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y133_IOB_X0Y133_IBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_IPAD),
.O(LIOB33_X0Y133_IOB_X0Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y133_IOB_X0Y134_IBUF (
.I(LIOB33_X0Y133_IOB_X0Y134_IPAD),
.O(LIOB33_X0Y133_IOB_X0Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y135_IOB_X0Y135_IBUF (
.I(LIOB33_X0Y135_IOB_X0Y135_IPAD),
.O(LIOB33_X0Y135_IOB_X0Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y135_IOB_X0Y136_IBUF (
.I(LIOB33_X0Y135_IOB_X0Y136_IPAD),
.O(LIOB33_X0Y135_IOB_X0Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(LIOB33_X0Y137_IOB_X0Y137_IPAD),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y137_IOB_X0Y138_IBUF (
.I(LIOB33_X0Y137_IOB_X0Y138_IPAD),
.O(LIOB33_X0Y137_IOB_X0Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y139_IOB_X0Y139_IBUF (
.I(LIOB33_X0Y139_IOB_X0Y139_IPAD),
.O(LIOB33_X0Y139_IOB_X0Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y139_IOB_X0Y140_IBUF (
.I(LIOB33_X0Y139_IOB_X0Y140_IPAD),
.O(LIOB33_X0Y139_IOB_X0Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y141_IOB_X0Y141_IBUF (
.I(LIOB33_X0Y141_IOB_X0Y141_IPAD),
.O(LIOB33_X0Y141_IOB_X0Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y141_IOB_X0Y142_IBUF (
.I(LIOB33_X0Y141_IOB_X0Y142_IPAD),
.O(LIOB33_X0Y141_IOB_X0Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y143_IOB_X0Y143_IBUF (
.I(LIOB33_X0Y143_IOB_X0Y143_IPAD),
.O(LIOB33_X0Y143_IOB_X0Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y145_IOB_X0Y145_IBUF (
.I(LIOB33_X0Y145_IOB_X0Y145_IPAD),
.O(LIOB33_X0Y145_IOB_X0Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y145_IOB_X0Y146_IBUF (
.I(LIOB33_X0Y145_IOB_X0Y146_IPAD),
.O(LIOB33_X0Y145_IOB_X0Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y147_IOB_X0Y147_IBUF (
.I(LIOB33_X0Y147_IOB_X0Y147_IPAD),
.O(LIOB33_X0Y147_IOB_X0Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y147_IOB_X0Y148_IBUF (
.I(LIOB33_X0Y147_IOB_X0Y148_IPAD),
.O(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y151_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y151_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y152_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y152_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y153_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y153_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y154_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y154_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y155_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y155_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y156_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y156_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y157_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y157_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y158_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y158_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y159_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y159_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y160_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y160_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y160_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y161_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y161_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y161_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y162_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y162_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y162_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y163_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y163_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y163_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y164_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y164_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y164_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y165_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y165_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y165_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y166_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y166_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y166_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y167_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y167_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y167_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y168_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y168_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y168_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y169_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y169_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y169_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y170_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y170_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y170_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y171_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y171_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y171_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y172_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y172_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y172_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y173_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y173_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y173_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y174_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y174_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y174_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y175_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y175_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y175_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y176_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y176_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y176_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y177_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y177_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y177_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y178_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y178_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y178_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y179_IOB_X0Y179_IBUF (
.I(LIOB33_X0Y179_IOB_X0Y179_IPAD),
.O(LIOB33_X0Y179_IOB_X0Y179_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y179_IOB_X0Y180_IBUF (
.I(LIOB33_X0Y179_IOB_X0Y180_IPAD),
.O(LIOB33_X0Y179_IOB_X0Y180_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y181_IOB_X0Y181_IBUF (
.I(LIOB33_X0Y181_IOB_X0Y181_IPAD),
.O(LIOB33_X0Y181_IOB_X0Y181_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y181_IOB_X0Y182_IBUF (
.I(LIOB33_X0Y181_IOB_X0Y182_IPAD),
.O(LIOB33_X0Y181_IOB_X0Y182_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y183_IOB_X0Y183_IBUF (
.I(LIOB33_X0Y183_IOB_X0Y183_IPAD),
.O(LIOB33_X0Y183_IOB_X0Y183_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y183_IOB_X0Y184_IBUF (
.I(LIOB33_X0Y183_IOB_X0Y184_IPAD),
.O(LIOB33_X0Y183_IOB_X0Y184_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y185_IOB_X0Y185_IBUF (
.I(LIOB33_X0Y185_IOB_X0Y185_IPAD),
.O(LIOB33_X0Y185_IOB_X0Y185_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y185_IOB_X0Y186_IBUF (
.I(LIOB33_X0Y185_IOB_X0Y186_IPAD),
.O(LIOB33_X0Y185_IOB_X0Y186_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y187_IOB_X0Y187_IBUF (
.I(LIOB33_X0Y187_IOB_X0Y187_IPAD),
.O(LIOB33_X0Y187_IOB_X0Y187_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y187_IOB_X0Y188_IBUF (
.I(LIOB33_X0Y187_IOB_X0Y188_IPAD),
.O(LIOB33_X0Y187_IOB_X0Y188_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y189_IOB_X0Y189_IBUF (
.I(LIOB33_X0Y189_IOB_X0Y189_IPAD),
.O(LIOB33_X0Y189_IOB_X0Y189_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y189_IOB_X0Y190_IBUF (
.I(LIOB33_X0Y189_IOB_X0Y190_IPAD),
.O(LIOB33_X0Y189_IOB_X0Y190_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y191_IOB_X0Y191_IBUF (
.I(LIOB33_X0Y191_IOB_X0Y191_IPAD),
.O(LIOB33_X0Y191_IOB_X0Y191_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y191_IOB_X0Y192_IBUF (
.I(LIOB33_X0Y191_IOB_X0Y192_IPAD),
.O(LIOB33_X0Y191_IOB_X0Y192_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y193_IOB_X0Y193_IBUF (
.I(LIOB33_X0Y193_IOB_X0Y193_IPAD),
.O(LIOB33_X0Y193_IOB_X0Y193_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y193_IOB_X0Y194_IBUF (
.I(LIOB33_X0Y193_IOB_X0Y194_IPAD),
.O(LIOB33_X0Y193_IOB_X0Y194_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y195_IOB_X0Y195_IBUF (
.I(LIOB33_X0Y195_IOB_X0Y195_IPAD),
.O(LIOB33_X0Y195_IOB_X0Y195_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y195_IOB_X0Y196_IBUF (
.I(LIOB33_X0Y195_IOB_X0Y196_IPAD),
.O(LIOB33_X0Y195_IOB_X0Y196_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y197_IOB_X0Y197_IBUF (
.I(LIOB33_X0Y197_IOB_X0Y197_IPAD),
.O(LIOB33_X0Y197_IOB_X0Y197_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y197_IOB_X0Y198_IBUF (
.I(LIOB33_X0Y197_IOB_X0Y198_IPAD),
.O(LIOB33_X0Y197_IOB_X0Y198_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y201_IOB_X0Y201_IBUF (
.I(LIOB33_X0Y201_IOB_X0Y201_IPAD),
.O(LIOB33_X0Y201_IOB_X0Y201_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y201_IOB_X0Y202_IBUF (
.I(LIOB33_X0Y201_IOB_X0Y202_IPAD),
.O(LIOB33_X0Y201_IOB_X0Y202_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y203_IOB_X0Y203_IBUF (
.I(LIOB33_X0Y203_IOB_X0Y203_IPAD),
.O(LIOB33_X0Y203_IOB_X0Y203_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y203_IOB_X0Y204_IBUF (
.I(LIOB33_X0Y203_IOB_X0Y204_IPAD),
.O(LIOB33_X0Y203_IOB_X0Y204_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y205_IOB_X0Y205_IBUF (
.I(LIOB33_X0Y205_IOB_X0Y205_IPAD),
.O(LIOB33_X0Y205_IOB_X0Y205_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y205_IOB_X0Y206_IBUF (
.I(LIOB33_X0Y205_IOB_X0Y206_IPAD),
.O(LIOB33_X0Y205_IOB_X0Y206_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y207_IOB_X0Y207_IBUF (
.I(LIOB33_X0Y207_IOB_X0Y207_IPAD),
.O(LIOB33_X0Y207_IOB_X0Y207_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y207_IOB_X0Y208_IBUF (
.I(LIOB33_X0Y207_IOB_X0Y208_IPAD),
.O(LIOB33_X0Y207_IOB_X0Y208_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y209_IOB_X0Y209_IBUF (
.I(LIOB33_X0Y209_IOB_X0Y209_IPAD),
.O(LIOB33_X0Y209_IOB_X0Y209_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y209_IOB_X0Y210_IBUF (
.I(LIOB33_X0Y209_IOB_X0Y210_IPAD),
.O(LIOB33_X0Y209_IOB_X0Y210_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y211_IOB_X0Y211_IBUF (
.I(LIOB33_X0Y211_IOB_X0Y211_IPAD),
.O(LIOB33_X0Y211_IOB_X0Y211_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y211_IOB_X0Y212_IBUF (
.I(LIOB33_X0Y211_IOB_X0Y212_IPAD),
.O(LIOB33_X0Y211_IOB_X0Y212_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y213_IOB_X0Y213_IBUF (
.I(LIOB33_X0Y213_IOB_X0Y213_IPAD),
.O(LIOB33_X0Y213_IOB_X0Y213_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y213_IOB_X0Y214_IBUF (
.I(LIOB33_X0Y213_IOB_X0Y214_IPAD),
.O(LIOB33_X0Y213_IOB_X0Y214_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y215_IOB_X0Y215_IBUF (
.I(LIOB33_X0Y215_IOB_X0Y215_IPAD),
.O(LIOB33_X0Y215_IOB_X0Y215_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y215_IOB_X0Y216_IBUF (
.I(LIOB33_X0Y215_IOB_X0Y216_IPAD),
.O(LIOB33_X0Y215_IOB_X0Y216_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y217_IOB_X0Y217_IBUF (
.I(LIOB33_X0Y217_IOB_X0Y217_IPAD),
.O(LIOB33_X0Y217_IOB_X0Y217_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y217_IOB_X0Y218_IBUF (
.I(LIOB33_X0Y217_IOB_X0Y218_IPAD),
.O(LIOB33_X0Y217_IOB_X0Y218_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y219_IOB_X0Y219_IBUF (
.I(LIOB33_X0Y219_IOB_X0Y219_IPAD),
.O(LIOB33_X0Y219_IOB_X0Y219_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y219_IOB_X0Y220_IBUF (
.I(LIOB33_X0Y219_IOB_X0Y220_IPAD),
.O(LIOB33_X0Y219_IOB_X0Y220_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y221_IOB_X0Y221_IBUF (
.I(LIOB33_X0Y221_IOB_X0Y221_IPAD),
.O(LIOB33_X0Y221_IOB_X0Y221_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y221_IOB_X0Y222_IBUF (
.I(LIOB33_X0Y221_IOB_X0Y222_IPAD),
.O(LIOB33_X0Y221_IOB_X0Y222_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y223_IOB_X0Y223_IBUF (
.I(LIOB33_X0Y223_IOB_X0Y223_IPAD),
.O(LIOB33_X0Y223_IOB_X0Y223_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y223_IOB_X0Y224_IBUF (
.I(LIOB33_X0Y223_IOB_X0Y224_IPAD),
.O(LIOB33_X0Y223_IOB_X0Y224_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y225_IOB_X0Y225_IBUF (
.I(LIOB33_X0Y225_IOB_X0Y225_IPAD),
.O(LIOB33_X0Y225_IOB_X0Y225_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y225_IOB_X0Y226_IBUF (
.I(LIOB33_X0Y225_IOB_X0Y226_IPAD),
.O(LIOB33_X0Y225_IOB_X0Y226_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y227_IOB_X0Y227_IBUF (
.I(LIOB33_X0Y227_IOB_X0Y227_IPAD),
.O(LIOB33_X0Y227_IOB_X0Y227_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y227_IOB_X0Y228_IBUF (
.I(LIOB33_X0Y227_IOB_X0Y228_IPAD),
.O(LIOB33_X0Y227_IOB_X0Y228_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y229_IOB_X0Y229_IBUF (
.I(LIOB33_X0Y229_IOB_X0Y229_IPAD),
.O(LIOB33_X0Y229_IOB_X0Y229_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y229_IOB_X0Y230_IBUF (
.I(LIOB33_X0Y229_IOB_X0Y230_IPAD),
.O(LIOB33_X0Y229_IOB_X0Y230_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y231_IOB_X0Y231_IBUF (
.I(LIOB33_X0Y231_IOB_X0Y231_IPAD),
.O(LIOB33_X0Y231_IOB_X0Y231_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y231_IOB_X0Y232_IBUF (
.I(LIOB33_X0Y231_IOB_X0Y232_IPAD),
.O(LIOB33_X0Y231_IOB_X0Y232_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y233_IOB_X0Y233_IBUF (
.I(LIOB33_X0Y233_IOB_X0Y233_IPAD),
.O(LIOB33_X0Y233_IOB_X0Y233_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y233_IOB_X0Y234_IBUF (
.I(LIOB33_X0Y233_IOB_X0Y234_IPAD),
.O(LIOB33_X0Y233_IOB_X0Y234_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y235_IOB_X0Y235_IBUF (
.I(LIOB33_X0Y235_IOB_X0Y235_IPAD),
.O(LIOB33_X0Y235_IOB_X0Y235_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y235_IOB_X0Y236_IBUF (
.I(LIOB33_X0Y235_IOB_X0Y236_IPAD),
.O(LIOB33_X0Y235_IOB_X0Y236_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y237_IOB_X0Y237_IBUF (
.I(LIOB33_X0Y237_IOB_X0Y237_IPAD),
.O(LIOB33_X0Y237_IOB_X0Y237_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y237_IOB_X0Y238_IBUF (
.I(LIOB33_X0Y237_IOB_X0Y238_IPAD),
.O(LIOB33_X0Y237_IOB_X0Y238_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y239_IOB_X0Y239_IBUF (
.I(LIOB33_X0Y239_IOB_X0Y239_IPAD),
.O(LIOB33_X0Y239_IOB_X0Y239_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y239_IOB_X0Y240_IBUF (
.I(LIOB33_X0Y239_IOB_X0Y240_IPAD),
.O(LIOB33_X0Y239_IOB_X0Y240_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y241_IOB_X0Y241_IBUF (
.I(LIOB33_X0Y241_IOB_X0Y241_IPAD),
.O(LIOB33_X0Y241_IOB_X0Y241_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y241_IOB_X0Y242_IBUF (
.I(LIOB33_X0Y241_IOB_X0Y242_IPAD),
.O(LIOB33_X0Y241_IOB_X0Y242_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y243_IOB_X0Y243_IBUF (
.I(LIOB33_X0Y243_IOB_X0Y243_IPAD),
.O(LIOB33_X0Y243_IOB_X0Y243_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y0_IOB_X0Y0_IBUF (
.I(LIOB33_SING_X0Y0_IOB_X0Y0_IPAD),
.O(LIOB33_SING_X0Y0_IOB_X0Y0_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y99_IOB_X0Y99_IBUF (
.I(LIOB33_SING_X0Y99_IOB_X0Y99_IPAD),
.O(LIOB33_SING_X0Y99_IOB_X0Y99_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y149_IOB_X0Y149_IBUF (
.I(LIOB33_SING_X0Y149_IOB_X0Y149_IPAD),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y150_IOB_X0Y150_IBUF (
.I(LIOB33_SING_X0Y150_IOB_X0Y150_IPAD),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y199_IOB_X0Y199_IBUF (
.I(LIOB33_SING_X0Y199_IOB_X0Y199_IPAD),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y200_IOB_X0Y200_IBUF (
.I(LIOB33_SING_X0Y200_IOB_X0Y200_IPAD),
.O(LIOB33_SING_X0Y200_IOB_X0Y200_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y51_IOB_X1Y51_OBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_I),
.O(RIOB33_X105Y51_IOB_X1Y51_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y51_IOB_X1Y52_OBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_I),
.O(RIOB33_X105Y51_IOB_X1Y52_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y53_IOB_X1Y53_OBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_I),
.O(RIOB33_X105Y53_IOB_X1Y53_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y53_IOB_X1Y54_OBUF (
.I(LIOB33_X0Y79_IOB_X0Y80_I),
.O(RIOB33_X105Y53_IOB_X1Y54_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y55_IOB_X1Y55_OBUF (
.I(CLBLL_L_X2Y103_SLICE_X1Y103_AO6),
.O(RIOB33_X105Y55_IOB_X1Y55_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y55_IOB_X1Y56_OBUF (
.I(CLBLL_L_X2Y104_SLICE_X0Y104_AO6),
.O(RIOB33_X105Y55_IOB_X1Y56_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y57_IOB_X1Y57_OBUF (
.I(CLBLL_L_X2Y210_SLICE_X0Y210_AO6),
.O(RIOB33_X105Y57_IOB_X1Y57_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y57_IOB_X1Y58_OBUF (
.I(LIOB33_X0Y81_IOB_X0Y82_I),
.O(RIOB33_X105Y57_IOB_X1Y58_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y59_IOB_X1Y59_OBUF (
.I(LIOB33_X0Y83_IOB_X0Y83_I),
.O(RIOB33_X105Y59_IOB_X1Y59_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y59_IOB_X1Y60_OBUF (
.I(LIOB33_X0Y83_IOB_X0Y84_I),
.O(RIOB33_X105Y59_IOB_X1Y60_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y61_IOB_X1Y61_OBUF (
.I(LIOB33_X0Y85_IOB_X0Y85_I),
.O(RIOB33_X105Y61_IOB_X1Y61_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y61_IOB_X1Y62_OBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_I),
.O(RIOB33_X105Y61_IOB_X1Y62_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y63_OBUF (
.I(LIOB33_X0Y85_IOB_X0Y86_I),
.O(RIOB33_X105Y63_IOB_X1Y63_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y64_OBUF (
.I(LIOB33_X0Y87_IOB_X0Y87_I),
.O(RIOB33_X105Y63_IOB_X1Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y65_OBUF (
.I(LIOB33_X0Y87_IOB_X0Y88_I),
.O(RIOB33_X105Y65_IOB_X1Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y66_OBUF (
.I(LIOB33_X0Y89_IOB_X0Y90_I),
.O(RIOB33_X105Y65_IOB_X1Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y67_OBUF (
.I(LIOB33_X0Y91_IOB_X0Y91_I),
.O(RIOB33_X105Y67_IOB_X1Y67_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y68_OBUF (
.I(LIOB33_X0Y91_IOB_X0Y92_I),
.O(RIOB33_X105Y67_IOB_X1Y68_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y69_OBUF (
.I(LIOB33_X0Y93_IOB_X0Y93_I),
.O(RIOB33_X105Y69_IOB_X1Y69_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y70_OBUF (
.I(LIOB33_X0Y93_IOB_X0Y94_I),
.O(RIOB33_X105Y69_IOB_X1Y70_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y71_OBUF (
.I(LIOB33_X0Y95_IOB_X0Y95_I),
.O(RIOB33_X105Y71_IOB_X1Y71_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y72_OBUF (
.I(CLBLL_L_X2Y189_SLICE_X0Y189_AO6),
.O(RIOB33_X105Y71_IOB_X1Y72_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y73_OBUF (
.I(LIOB33_X0Y95_IOB_X0Y96_I),
.O(RIOB33_X105Y73_IOB_X1Y73_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y74_OBUF (
.I(CLBLM_L_X44Y158_SLICE_X66Y158_BO6),
.O(RIOB33_X105Y73_IOB_X1Y74_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y75_OBUF (
.I(CLBLM_L_X44Y152_SLICE_X66Y152_AO6),
.O(RIOB33_X105Y75_IOB_X1Y75_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y76_OBUF (
.I(LIOB33_X0Y97_IOB_X0Y97_I),
.O(RIOB33_X105Y75_IOB_X1Y76_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y77_IOB_X1Y77_OBUF (
.I(LIOB33_X0Y97_IOB_X0Y98_I),
.O(RIOB33_X105Y77_IOB_X1Y77_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y77_IOB_X1Y78_OBUF (
.I(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.O(RIOB33_X105Y77_IOB_X1Y78_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y79_OBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_I),
.O(RIOB33_X105Y79_IOB_X1Y79_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y80_OBUF (
.I(CLBLL_L_X2Y208_SLICE_X0Y208_AO6),
.O(RIOB33_X105Y79_IOB_X1Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y81_OBUF (
.I(CLBLL_L_X2Y210_SLICE_X0Y210_AO6),
.O(RIOB33_X105Y81_IOB_X1Y81_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y82_OBUF (
.I(CLBLL_L_X2Y193_SLICE_X0Y193_AO6),
.O(RIOB33_X105Y81_IOB_X1Y82_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y83_OBUF (
.I(CLBLL_L_X2Y189_SLICE_X1Y189_AO6),
.O(RIOB33_X105Y83_IOB_X1Y83_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y84_OBUF (
.I(CLBLL_L_X2Y187_SLICE_X0Y187_AO6),
.O(RIOB33_X105Y83_IOB_X1Y84_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y85_OBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_I),
.O(RIOB33_X105Y85_IOB_X1Y85_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y86_OBUF (
.I(CLBLL_L_X2Y194_SLICE_X0Y194_AO6),
.O(RIOB33_X105Y85_IOB_X1Y86_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y87_OBUF (
.I(CLBLL_L_X2Y192_SLICE_X0Y192_AO6),
.O(RIOB33_X105Y87_IOB_X1Y87_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y88_OBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_I),
.O(RIOB33_X105Y87_IOB_X1Y88_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y89_OBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_I),
.O(RIOB33_X105Y89_IOB_X1Y89_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y90_OBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_I),
.O(RIOB33_X105Y89_IOB_X1Y90_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y91_OBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_I),
.O(RIOB33_X105Y91_IOB_X1Y91_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y92_OBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_I),
.O(RIOB33_X105Y91_IOB_X1Y92_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y93_IOB_X1Y93_OBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_I),
.O(RIOB33_X105Y93_IOB_X1Y93_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y93_IOB_X1Y94_OBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_I),
.O(RIOB33_X105Y93_IOB_X1Y94_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y95_IOB_X1Y95_OBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_I),
.O(RIOB33_X105Y95_IOB_X1Y95_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y95_IOB_X1Y96_OBUF (
.I(LIOB33_X0Y119_IOB_X0Y120_I),
.O(RIOB33_X105Y95_IOB_X1Y96_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y97_IOB_X1Y97_OBUF (
.I(LIOB33_X0Y121_IOB_X0Y121_I),
.O(RIOB33_X105Y97_IOB_X1Y97_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y97_IOB_X1Y98_OBUF (
.I(LIOB33_X0Y121_IOB_X0Y122_I),
.O(RIOB33_X105Y97_IOB_X1Y98_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y101_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_I),
.O(RIOB33_X105Y101_IOB_X1Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y102_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(RIOB33_X105Y101_IOB_X1Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y103_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_X105Y103_IOB_X1Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y104_OBUF (
.I(CLBLL_L_X2Y103_SLICE_X0Y103_AO6),
.O(RIOB33_X105Y103_IOB_X1Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y105_OBUF (
.I(CLBLL_L_X2Y189_SLICE_X1Y189_AO6),
.O(RIOB33_X105Y105_IOB_X1Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y106_OBUF (
.I(LIOB33_X0Y81_IOB_X0Y81_I),
.O(RIOB33_X105Y105_IOB_X1Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y107_OBUF (
.I(LIOB33_X0Y201_IOB_X0Y201_I),
.O(RIOB33_X105Y107_IOB_X1Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y108_OBUF (
.I(LIOB33_X0Y201_IOB_X0Y202_I),
.O(RIOB33_X105Y107_IOB_X1Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y109_OBUF (
.I(LIOB33_X0Y203_IOB_X0Y203_I),
.O(RIOB33_X105Y109_IOB_X1Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y110_OBUF (
.I(LIOB33_X0Y203_IOB_X0Y204_I),
.O(RIOB33_X105Y109_IOB_X1Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y111_OBUF (
.I(LIOB33_X0Y205_IOB_X0Y205_I),
.O(RIOB33_X105Y111_IOB_X1Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y112_OBUF (
.I(CLBLL_L_X2Y192_SLICE_X0Y192_BO6),
.O(RIOB33_X105Y111_IOB_X1Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y113_OBUF (
.I(CLBLL_L_X2Y192_SLICE_X0Y192_BO6),
.O(RIOB33_X105Y113_IOB_X1Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y114_OBUF (
.I(CLBLL_L_X2Y193_SLICE_X0Y193_BO6),
.O(RIOB33_X105Y113_IOB_X1Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y115_OBUF (
.I(CLBLL_L_X2Y193_SLICE_X0Y193_BO6),
.O(RIOB33_X105Y115_IOB_X1Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y116_OBUF (
.I(CLBLL_L_X2Y192_SLICE_X0Y192_CO6),
.O(RIOB33_X105Y115_IOB_X1Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y117_OBUF (
.I(CLBLL_L_X2Y150_SLICE_X0Y150_CO6),
.O(RIOB33_X105Y117_IOB_X1Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y118_OBUF (
.I(CLBLL_L_X2Y150_SLICE_X0Y150_CO6),
.O(RIOB33_X105Y117_IOB_X1Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y119_OBUF (
.I(CLBLL_L_X2Y138_SLICE_X0Y138_AO6),
.O(RIOB33_X105Y119_IOB_X1Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y120_OBUF (
.I(CLBLM_R_X67Y130_SLICE_X100Y130_AO6),
.O(RIOB33_X105Y119_IOB_X1Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y121_OBUF (
.I(CLBLL_L_X2Y154_SLICE_X0Y154_AO6),
.O(RIOB33_X105Y121_IOB_X1Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y122_OBUF (
.I(CLBLL_L_X2Y145_SLICE_X0Y145_AO6),
.O(RIOB33_X105Y121_IOB_X1Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y123_OBUF (
.I(CLBLL_L_X2Y142_SLICE_X0Y142_CO6),
.O(RIOB33_X105Y123_IOB_X1Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y124_OBUF (
.I(CLBLL_L_X2Y142_SLICE_X0Y142_CO6),
.O(RIOB33_X105Y123_IOB_X1Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y125_OBUF (
.I(1'b1),
.O(RIOB33_X105Y125_IOB_X1Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y126_OBUF (
.I(CLBLL_L_X2Y134_SLICE_X0Y134_AO6),
.O(RIOB33_X105Y125_IOB_X1Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(CLBLL_L_X2Y151_SLICE_X0Y151_BO6),
.O(RIOB33_X105Y127_IOB_X1Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y128_OBUF (
.I(CLBLL_L_X2Y151_SLICE_X0Y151_BO6),
.O(RIOB33_X105Y127_IOB_X1Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(CLBLL_L_X2Y151_SLICE_X0Y151_CO6),
.O(RIOB33_X105Y129_IOB_X1Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(CLBLL_L_X2Y148_SLICE_X0Y148_DO6),
.O(RIOB33_X105Y129_IOB_X1Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(1'b0),
.O(RIOB33_X105Y131_IOB_X1Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(CLBLM_R_X59Y133_SLICE_X88Y133_AO6),
.O(RIOB33_X105Y131_IOB_X1Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(CLBLM_R_X59Y133_SLICE_X88Y133_AO6),
.O(RIOB33_X105Y133_IOB_X1Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_I),
.O(RIOB33_X105Y133_IOB_X1Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_I),
.O(RIOB33_X105Y135_IOB_X1Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y136_OBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_I),
.O(RIOB33_X105Y135_IOB_X1Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y137_OBUF (
.I(LIOB33_X0Y135_IOB_X0Y135_I),
.O(RIOB33_X105Y137_IOB_X1Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y138_OBUF (
.I(LIOB33_X0Y135_IOB_X0Y135_I),
.O(RIOB33_X105Y137_IOB_X1Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y139_OBUF (
.I(LIOB33_X0Y155_IOB_X0Y155_I),
.O(RIOB33_X105Y139_IOB_X1Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y140_OBUF (
.I(LIOB33_X0Y183_IOB_X0Y184_I),
.O(RIOB33_X105Y139_IOB_X1Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y141_OBUF (
.I(LIOB33_X0Y9_IOB_X0Y10_I),
.O(RIOB33_X105Y141_IOB_X1Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y142_OBUF (
.I(LIOB33_X0Y229_IOB_X0Y230_I),
.O(RIOB33_X105Y141_IOB_X1Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y143_OBUF (
.I(LIOB33_X0Y217_IOB_X0Y217_I),
.O(RIOB33_X105Y143_IOB_X1Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y144_OBUF (
.I(LIOB33_X0Y1_IOB_X0Y1_I),
.O(RIOB33_X105Y143_IOB_X1Y144_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y145_OBUF (
.I(LIOB33_X0Y195_IOB_X0Y195_I),
.O(RIOB33_X105Y145_IOB_X1Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y146_OBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_I),
.O(RIOB33_X105Y145_IOB_X1Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y147_OBUF (
.I(CLBLL_L_X2Y149_SLICE_X0Y149_AO5),
.O(RIOB33_X105Y147_IOB_X1Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y148_OBUF (
.I(CLBLL_L_X2Y147_SLICE_X0Y147_BO6),
.O(RIOB33_X105Y147_IOB_X1Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y151_IOB_X1Y151_IBUF (
.I(RIOB33_X105Y151_IOB_X1Y151_IPAD),
.O(RIOB33_X105Y151_IOB_X1Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y151_IOB_X1Y152_IBUF (
.I(RIOB33_X105Y151_IOB_X1Y152_IPAD),
.O(RIOB33_X105Y151_IOB_X1Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y153_IOB_X1Y153_IBUF (
.I(RIOB33_X105Y153_IOB_X1Y153_IPAD),
.O(RIOB33_X105Y153_IOB_X1Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y153_IOB_X1Y154_IBUF (
.I(RIOB33_X105Y153_IOB_X1Y154_IPAD),
.O(RIOB33_X105Y153_IOB_X1Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y155_IOB_X1Y155_IBUF (
.I(RIOB33_X105Y155_IOB_X1Y155_IPAD),
.O(RIOB33_X105Y155_IOB_X1Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y155_IOB_X1Y156_IBUF (
.I(RIOB33_X105Y155_IOB_X1Y156_IPAD),
.O(RIOB33_X105Y155_IOB_X1Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y157_IOB_X1Y157_IBUF (
.I(RIOB33_X105Y157_IOB_X1Y157_IPAD),
.O(RIOB33_X105Y157_IOB_X1Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y157_IOB_X1Y158_IBUF (
.I(RIOB33_X105Y157_IOB_X1Y158_IPAD),
.O(RIOB33_X105Y157_IOB_X1Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y159_IOB_X1Y159_IBUF (
.I(RIOB33_X105Y159_IOB_X1Y159_IPAD),
.O(RIOB33_X105Y159_IOB_X1Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_R_X59Y159_SLICE_X88Y159_AO6),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X44Y158_SLICE_X66Y158_BO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X44Y158_SLICE_X66Y158_AO5),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X44Y158_SLICE_X66Y158_AO6),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_R_X47Y158_SLICE_X72Y158_AO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(LIOB33_X0Y19_IOB_X0Y19_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(CLBLM_R_X47Y158_SLICE_X72Y158_AO5),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_X0Y19_IOB_X0Y20_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(LIOB33_X0Y21_IOB_X0Y21_I),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(LIOB33_X0Y21_IOB_X0Y22_I),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(LIOB33_X0Y23_IOB_X0Y23_I),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(LIOB33_X0Y23_IOB_X0Y24_I),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(LIOB33_X0Y25_IOB_X0Y25_I),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(LIOB33_X0Y27_IOB_X0Y27_I),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(LIOB33_X0Y27_IOB_X0Y28_I),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_I),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_I),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X44Y152_SLICE_X66Y152_AO5),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLL_L_X2Y193_SLICE_X0Y193_AO6),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(LIOB33_X0Y155_IOB_X0Y155_I),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(LIOB33_X0Y155_IOB_X0Y155_I),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y50_IOB_X1Y50_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_SING_X105Y50_IOB_X1Y50_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y99_IOB_X1Y99_OBUF (
.I(LIOB33_SING_X0Y200_IOB_X0Y200_I),
.O(RIOB33_SING_X105Y99_IOB_X1Y99_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y100_IOB_X1Y100_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y149_IOB_X1Y149_OBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_I),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y150_IOB_X1Y150_IBUF (
.I(RIOB33_SING_X105Y150_IOB_X1Y150_IPAD),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(LIOB33_X0Y241_IOB_X0Y242_I),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A = CLBLL_L_X2Y102_SLICE_X0Y102_AO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B = CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C = CLBLL_L_X2Y102_SLICE_X0Y102_CO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D = CLBLL_L_X2Y102_SLICE_X0Y102_DO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A = CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B = CLBLL_L_X2Y102_SLICE_X1Y102_BO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C = CLBLL_L_X2Y102_SLICE_X1Y102_CO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D = CLBLL_L_X2Y102_SLICE_X1Y102_DO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B = CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C = CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D = CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A = CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D = CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A = CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C = CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D = CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D = CLBLL_L_X2Y130_SLICE_X0Y130_DO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A = CLBLL_L_X2Y130_SLICE_X1Y130_AO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B = CLBLL_L_X2Y130_SLICE_X1Y130_BO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C = CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D = CLBLL_L_X2Y130_SLICE_X1Y130_DO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B = CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C = CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D = CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A = CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B = CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C = CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D = CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A = CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B = CLBLL_L_X2Y134_SLICE_X0Y134_BO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C = CLBLL_L_X2Y134_SLICE_X0Y134_CO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D = CLBLL_L_X2Y134_SLICE_X0Y134_DO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A = CLBLL_L_X2Y134_SLICE_X1Y134_AO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B = CLBLL_L_X2Y134_SLICE_X1Y134_BO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C = CLBLL_L_X2Y134_SLICE_X1Y134_CO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D = CLBLL_L_X2Y134_SLICE_X1Y134_DO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B = CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C = CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D = CLBLL_L_X2Y138_SLICE_X0Y138_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A = CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B = CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C = CLBLL_L_X2Y138_SLICE_X1Y138_CO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D = CLBLL_L_X2Y138_SLICE_X1Y138_DO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A = CLBLL_L_X2Y142_SLICE_X0Y142_AO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B = CLBLL_L_X2Y142_SLICE_X0Y142_BO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C = CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D = CLBLL_L_X2Y142_SLICE_X0Y142_DO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A = CLBLL_L_X2Y142_SLICE_X1Y142_AO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B = CLBLL_L_X2Y142_SLICE_X1Y142_BO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C = CLBLL_L_X2Y142_SLICE_X1Y142_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D = CLBLL_L_X2Y142_SLICE_X1Y142_DO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A = CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B = CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C = CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D = CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A = CLBLL_L_X2Y145_SLICE_X1Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B = CLBLL_L_X2Y145_SLICE_X1Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C = CLBLL_L_X2Y145_SLICE_X1Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D = CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B = CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C = CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D = CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C = CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D = CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A = CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B = CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C = CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D = CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D = CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A = CLBLL_L_X2Y149_SLICE_X0Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B = CLBLL_L_X2Y149_SLICE_X0Y149_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C = CLBLL_L_X2Y149_SLICE_X0Y149_CO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D = CLBLL_L_X2Y149_SLICE_X0Y149_DO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_AMUX = CLBLL_L_X2Y149_SLICE_X0Y149_AO5;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A = CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B = CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C = CLBLL_L_X2Y149_SLICE_X1Y149_CO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D = CLBLL_L_X2Y149_SLICE_X1Y149_DO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_AMUX = CLBLL_L_X2Y149_SLICE_X1Y149_AO5;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_BMUX = CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A = CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B = CLBLL_L_X2Y150_SLICE_X0Y150_BO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C = CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D = CLBLL_L_X2Y150_SLICE_X0Y150_DO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A = CLBLL_L_X2Y150_SLICE_X1Y150_AO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B = CLBLL_L_X2Y150_SLICE_X1Y150_BO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C = CLBLL_L_X2Y150_SLICE_X1Y150_CO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D = CLBLL_L_X2Y150_SLICE_X1Y150_DO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A = CLBLL_L_X2Y151_SLICE_X0Y151_AO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C = CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D = CLBLL_L_X2Y151_SLICE_X0Y151_DO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A = CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C = CLBLL_L_X2Y151_SLICE_X1Y151_CO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D = CLBLL_L_X2Y151_SLICE_X1Y151_DO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A = CLBLL_L_X2Y154_SLICE_X0Y154_AO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B = CLBLL_L_X2Y154_SLICE_X0Y154_BO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C = CLBLL_L_X2Y154_SLICE_X0Y154_CO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D = CLBLL_L_X2Y154_SLICE_X0Y154_DO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C = CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D = CLBLL_L_X2Y154_SLICE_X1Y154_DO6;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_A = CLBLL_L_X2Y165_SLICE_X0Y165_AO6;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_B = CLBLL_L_X2Y165_SLICE_X0Y165_BO6;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_C = CLBLL_L_X2Y165_SLICE_X0Y165_CO6;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_D = CLBLL_L_X2Y165_SLICE_X0Y165_DO6;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_A = CLBLL_L_X2Y165_SLICE_X1Y165_AO6;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_B = CLBLL_L_X2Y165_SLICE_X1Y165_BO6;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_C = CLBLL_L_X2Y165_SLICE_X1Y165_CO6;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_D = CLBLL_L_X2Y165_SLICE_X1Y165_DO6;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_A = CLBLL_L_X2Y170_SLICE_X0Y170_AO6;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_B = CLBLL_L_X2Y170_SLICE_X0Y170_BO6;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_C = CLBLL_L_X2Y170_SLICE_X0Y170_CO6;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_D = CLBLL_L_X2Y170_SLICE_X0Y170_DO6;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_A = CLBLL_L_X2Y170_SLICE_X1Y170_AO6;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_B = CLBLL_L_X2Y170_SLICE_X1Y170_BO6;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_C = CLBLL_L_X2Y170_SLICE_X1Y170_CO6;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_D = CLBLL_L_X2Y170_SLICE_X1Y170_DO6;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_A = CLBLL_L_X2Y187_SLICE_X0Y187_AO6;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_B = CLBLL_L_X2Y187_SLICE_X0Y187_BO6;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_C = CLBLL_L_X2Y187_SLICE_X0Y187_CO6;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_D = CLBLL_L_X2Y187_SLICE_X0Y187_DO6;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_AMUX = CLBLL_L_X2Y187_SLICE_X0Y187_AO5;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_A = CLBLL_L_X2Y187_SLICE_X1Y187_AO6;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_B = CLBLL_L_X2Y187_SLICE_X1Y187_BO6;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_C = CLBLL_L_X2Y187_SLICE_X1Y187_CO6;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_D = CLBLL_L_X2Y187_SLICE_X1Y187_DO6;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_A = CLBLL_L_X2Y189_SLICE_X0Y189_AO6;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_B = CLBLL_L_X2Y189_SLICE_X0Y189_BO6;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_C = CLBLL_L_X2Y189_SLICE_X0Y189_CO6;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_D = CLBLL_L_X2Y189_SLICE_X0Y189_DO6;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_A = CLBLL_L_X2Y189_SLICE_X1Y189_AO6;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_B = CLBLL_L_X2Y189_SLICE_X1Y189_BO6;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_C = CLBLL_L_X2Y189_SLICE_X1Y189_CO6;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_D = CLBLL_L_X2Y189_SLICE_X1Y189_DO6;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_A = CLBLL_L_X2Y192_SLICE_X0Y192_AO6;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_B = CLBLL_L_X2Y192_SLICE_X0Y192_BO6;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_C = CLBLL_L_X2Y192_SLICE_X0Y192_CO6;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_D = CLBLL_L_X2Y192_SLICE_X0Y192_DO6;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_A = CLBLL_L_X2Y192_SLICE_X1Y192_AO6;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_B = CLBLL_L_X2Y192_SLICE_X1Y192_BO6;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_C = CLBLL_L_X2Y192_SLICE_X1Y192_CO6;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_D = CLBLL_L_X2Y192_SLICE_X1Y192_DO6;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_A = CLBLL_L_X2Y193_SLICE_X0Y193_AO6;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_B = CLBLL_L_X2Y193_SLICE_X0Y193_BO6;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_C = CLBLL_L_X2Y193_SLICE_X0Y193_CO6;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_D = CLBLL_L_X2Y193_SLICE_X0Y193_DO6;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_A = CLBLL_L_X2Y193_SLICE_X1Y193_AO6;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_B = CLBLL_L_X2Y193_SLICE_X1Y193_BO6;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_C = CLBLL_L_X2Y193_SLICE_X1Y193_CO6;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_D = CLBLL_L_X2Y193_SLICE_X1Y193_DO6;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_A = CLBLL_L_X2Y194_SLICE_X0Y194_AO6;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_B = CLBLL_L_X2Y194_SLICE_X0Y194_BO6;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_C = CLBLL_L_X2Y194_SLICE_X0Y194_CO6;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_D = CLBLL_L_X2Y194_SLICE_X0Y194_DO6;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_A = CLBLL_L_X2Y194_SLICE_X1Y194_AO6;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_B = CLBLL_L_X2Y194_SLICE_X1Y194_BO6;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_C = CLBLL_L_X2Y194_SLICE_X1Y194_CO6;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_D = CLBLL_L_X2Y194_SLICE_X1Y194_DO6;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_A = CLBLL_L_X2Y208_SLICE_X0Y208_AO6;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_B = CLBLL_L_X2Y208_SLICE_X0Y208_BO6;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_C = CLBLL_L_X2Y208_SLICE_X0Y208_CO6;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_D = CLBLL_L_X2Y208_SLICE_X0Y208_DO6;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_A = CLBLL_L_X2Y208_SLICE_X1Y208_AO6;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_B = CLBLL_L_X2Y208_SLICE_X1Y208_BO6;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_C = CLBLL_L_X2Y208_SLICE_X1Y208_CO6;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_D = CLBLL_L_X2Y208_SLICE_X1Y208_DO6;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_A = CLBLL_L_X2Y210_SLICE_X0Y210_AO6;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_B = CLBLL_L_X2Y210_SLICE_X0Y210_BO6;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_C = CLBLL_L_X2Y210_SLICE_X0Y210_CO6;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_D = CLBLL_L_X2Y210_SLICE_X0Y210_DO6;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_A = CLBLL_L_X2Y210_SLICE_X1Y210_AO6;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_B = CLBLL_L_X2Y210_SLICE_X1Y210_BO6;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_C = CLBLL_L_X2Y210_SLICE_X1Y210_CO6;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_D = CLBLL_L_X2Y210_SLICE_X1Y210_DO6;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_A = CLBLM_L_X44Y152_SLICE_X66Y152_AO6;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_B = CLBLM_L_X44Y152_SLICE_X66Y152_BO6;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_C = CLBLM_L_X44Y152_SLICE_X66Y152_CO6;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_D = CLBLM_L_X44Y152_SLICE_X66Y152_DO6;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_AMUX = CLBLM_L_X44Y152_SLICE_X66Y152_AO5;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_A = CLBLM_L_X44Y152_SLICE_X67Y152_AO6;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_B = CLBLM_L_X44Y152_SLICE_X67Y152_BO6;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_C = CLBLM_L_X44Y152_SLICE_X67Y152_CO6;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_D = CLBLM_L_X44Y152_SLICE_X67Y152_DO6;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_A = CLBLM_L_X44Y158_SLICE_X66Y158_AO6;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_B = CLBLM_L_X44Y158_SLICE_X66Y158_BO6;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_C = CLBLM_L_X44Y158_SLICE_X66Y158_CO6;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_D = CLBLM_L_X44Y158_SLICE_X66Y158_DO6;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_AMUX = CLBLM_L_X44Y158_SLICE_X66Y158_AO5;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_BMUX = CLBLM_L_X44Y158_SLICE_X66Y158_BO5;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_A = CLBLM_L_X44Y158_SLICE_X67Y158_AO6;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_B = CLBLM_L_X44Y158_SLICE_X67Y158_BO6;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_C = CLBLM_L_X44Y158_SLICE_X67Y158_CO6;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_D = CLBLM_L_X44Y158_SLICE_X67Y158_DO6;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_A = CLBLM_R_X47Y145_SLICE_X72Y145_AO6;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_B = CLBLM_R_X47Y145_SLICE_X72Y145_BO6;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_C = CLBLM_R_X47Y145_SLICE_X72Y145_CO6;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_D = CLBLM_R_X47Y145_SLICE_X72Y145_DO6;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_A = CLBLM_R_X47Y145_SLICE_X73Y145_AO6;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_B = CLBLM_R_X47Y145_SLICE_X73Y145_BO6;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_C = CLBLM_R_X47Y145_SLICE_X73Y145_CO6;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_D = CLBLM_R_X47Y145_SLICE_X73Y145_DO6;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_A = CLBLM_R_X47Y158_SLICE_X72Y158_AO6;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_B = CLBLM_R_X47Y158_SLICE_X72Y158_BO6;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_C = CLBLM_R_X47Y158_SLICE_X72Y158_CO6;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_D = CLBLM_R_X47Y158_SLICE_X72Y158_DO6;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_AMUX = CLBLM_R_X47Y158_SLICE_X72Y158_AO5;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_A = CLBLM_R_X47Y158_SLICE_X73Y158_AO6;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_B = CLBLM_R_X47Y158_SLICE_X73Y158_BO6;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_C = CLBLM_R_X47Y158_SLICE_X73Y158_CO6;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_D = CLBLM_R_X47Y158_SLICE_X73Y158_DO6;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_A = CLBLM_R_X59Y133_SLICE_X88Y133_AO6;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_B = CLBLM_R_X59Y133_SLICE_X88Y133_BO6;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_C = CLBLM_R_X59Y133_SLICE_X88Y133_CO6;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_D = CLBLM_R_X59Y133_SLICE_X88Y133_DO6;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_A = CLBLM_R_X59Y133_SLICE_X89Y133_AO6;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_B = CLBLM_R_X59Y133_SLICE_X89Y133_BO6;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_C = CLBLM_R_X59Y133_SLICE_X89Y133_CO6;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_D = CLBLM_R_X59Y133_SLICE_X89Y133_DO6;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_A = CLBLM_R_X59Y159_SLICE_X88Y159_AO6;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_B = CLBLM_R_X59Y159_SLICE_X88Y159_BO6;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_C = CLBLM_R_X59Y159_SLICE_X88Y159_CO6;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_D = CLBLM_R_X59Y159_SLICE_X88Y159_DO6;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_A = CLBLM_R_X59Y159_SLICE_X89Y159_AO6;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_B = CLBLM_R_X59Y159_SLICE_X89Y159_BO6;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_C = CLBLM_R_X59Y159_SLICE_X89Y159_CO6;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_D = CLBLM_R_X59Y159_SLICE_X89Y159_DO6;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_A = CLBLM_R_X67Y130_SLICE_X100Y130_AO6;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_B = CLBLM_R_X67Y130_SLICE_X100Y130_BO6;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_C = CLBLM_R_X67Y130_SLICE_X100Y130_CO6;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_D = CLBLM_R_X67Y130_SLICE_X100Y130_DO6;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_A = CLBLM_R_X67Y130_SLICE_X101Y130_AO6;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_B = CLBLM_R_X67Y130_SLICE_X101Y130_BO6;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_C = CLBLM_R_X67Y130_SLICE_X101Y130_CO6;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_D = CLBLM_R_X67Y130_SLICE_X101Y130_DO6;
  assign LIOI3_X0Y1_ILOGIC_X0Y2_O = LIOB33_X0Y1_IOB_X0Y2_I;
  assign LIOI3_X0Y1_ILOGIC_X0Y1_O = LIOB33_X0Y1_IOB_X0Y1_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y4_O = LIOB33_X0Y3_IOB_X0Y4_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y3_O = LIOB33_X0Y3_IOB_X0Y3_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_O = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_O = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_O = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_O = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_O = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_O = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_O = LIOB33_X0Y15_IOB_X0Y16_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_O = LIOB33_X0Y15_IOB_X0Y15_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_O = LIOB33_X0Y17_IOB_X0Y18_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_O = LIOB33_X0Y17_IOB_X0Y17_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_O = LIOB33_X0Y21_IOB_X0Y22_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_O = LIOB33_X0Y21_IOB_X0Y21_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_O = LIOB33_X0Y23_IOB_X0Y24_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_O = LIOB33_X0Y23_IOB_X0Y23_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_O = LIOB33_X0Y25_IOB_X0Y26_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_O = LIOB33_X0Y25_IOB_X0Y25_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_O = LIOB33_X0Y27_IOB_X0Y28_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_O = LIOB33_X0Y27_IOB_X0Y27_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y80_O = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y84_O = LIOB33_X0Y83_IOB_X0Y84_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y83_O = LIOB33_X0Y83_IOB_X0Y83_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y86_O = LIOB33_X0Y85_IOB_X0Y86_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y85_O = LIOB33_X0Y85_IOB_X0Y85_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y90_O = LIOB33_X0Y89_IOB_X0Y90_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y89_O = LIOB33_X0Y89_IOB_X0Y89_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y92_O = LIOB33_X0Y91_IOB_X0Y92_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y91_O = LIOB33_X0Y91_IOB_X0Y91_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y96_O = LIOB33_X0Y95_IOB_X0Y96_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y95_O = LIOB33_X0Y95_IOB_X0Y95_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y98_O = LIOB33_X0Y97_IOB_X0Y98_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y97_O = LIOB33_X0Y97_IOB_X0Y97_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_O = LIOB33_X0Y129_IOB_X0Y130_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_O = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_O = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y136_O = LIOB33_X0Y135_IOB_X0Y136_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_O = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y140_O = LIOB33_X0Y139_IOB_X0Y140_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y139_O = LIOB33_X0Y139_IOB_X0Y139_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_O = LIOB33_X0Y141_IOB_X0Y142_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_O = LIOB33_X0Y141_IOB_X0Y141_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_O = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_O = LIOB33_X0Y145_IOB_X0Y145_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y148_O = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_O = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_O = LIOB33_X0Y151_IOB_X0Y151_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_O = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_O = LIOB33_X0Y153_IOB_X0Y153_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_O = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_O = LIOB33_X0Y155_IOB_X0Y155_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_O = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_O = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_O = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_O = LIOB33_X0Y161_IOB_X0Y161_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_O = LIOB33_X0Y165_IOB_X0Y166_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_O = LIOB33_X0Y165_IOB_X0Y165_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y168_O = LIOB33_X0Y167_IOB_X0Y168_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_O = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_O = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_O = LIOB33_X0Y173_IOB_X0Y173_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_O = LIOB33_X0Y175_IOB_X0Y175_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y178_O = LIOB33_X0Y177_IOB_X0Y178_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_O = LIOB33_X0Y177_IOB_X0Y177_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y180_O = LIOB33_X0Y179_IOB_X0Y180_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y179_O = LIOB33_X0Y179_IOB_X0Y179_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y184_O = LIOB33_X0Y183_IOB_X0Y184_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y183_O = LIOB33_X0Y183_IOB_X0Y183_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y186_O = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y185_O = LIOB33_X0Y185_IOB_X0Y185_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y190_O = LIOB33_X0Y189_IOB_X0Y190_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y189_O = LIOB33_X0Y189_IOB_X0Y189_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y192_O = LIOB33_X0Y191_IOB_X0Y192_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y191_O = LIOB33_X0Y191_IOB_X0Y191_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y196_O = LIOB33_X0Y195_IOB_X0Y196_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y195_O = LIOB33_X0Y195_IOB_X0Y195_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y198_O = LIOB33_X0Y197_IOB_X0Y198_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y197_O = LIOB33_X0Y197_IOB_X0Y197_I;
  assign LIOI3_X0Y201_ILOGIC_X0Y202_O = LIOB33_X0Y201_IOB_X0Y202_I;
  assign LIOI3_X0Y201_ILOGIC_X0Y201_O = LIOB33_X0Y201_IOB_X0Y201_I;
  assign LIOI3_X0Y203_ILOGIC_X0Y204_O = LIOB33_X0Y203_IOB_X0Y204_I;
  assign LIOI3_X0Y203_ILOGIC_X0Y203_O = LIOB33_X0Y203_IOB_X0Y203_I;
  assign LIOI3_X0Y205_ILOGIC_X0Y206_O = LIOB33_X0Y205_IOB_X0Y206_I;
  assign LIOI3_X0Y205_ILOGIC_X0Y205_O = LIOB33_X0Y205_IOB_X0Y205_I;
  assign LIOI3_X0Y209_ILOGIC_X0Y210_O = LIOB33_X0Y209_IOB_X0Y210_I;
  assign LIOI3_X0Y209_ILOGIC_X0Y209_O = LIOB33_X0Y209_IOB_X0Y209_I;
  assign LIOI3_X0Y211_ILOGIC_X0Y212_O = LIOB33_X0Y211_IOB_X0Y212_I;
  assign LIOI3_X0Y211_ILOGIC_X0Y211_O = LIOB33_X0Y211_IOB_X0Y211_I;
  assign LIOI3_X0Y215_ILOGIC_X0Y216_O = LIOB33_X0Y215_IOB_X0Y216_I;
  assign LIOI3_X0Y215_ILOGIC_X0Y215_O = LIOB33_X0Y215_IOB_X0Y215_I;
  assign LIOI3_X0Y217_ILOGIC_X0Y218_O = LIOB33_X0Y217_IOB_X0Y218_I;
  assign LIOI3_X0Y217_ILOGIC_X0Y217_O = LIOB33_X0Y217_IOB_X0Y217_I;
  assign LIOI3_X0Y221_ILOGIC_X0Y222_O = LIOB33_X0Y221_IOB_X0Y222_I;
  assign LIOI3_X0Y223_ILOGIC_X0Y224_O = LIOB33_X0Y223_IOB_X0Y224_I;
  assign LIOI3_X0Y223_ILOGIC_X0Y223_O = LIOB33_X0Y223_IOB_X0Y223_I;
  assign LIOI3_X0Y225_ILOGIC_X0Y226_O = LIOB33_X0Y225_IOB_X0Y226_I;
  assign LIOI3_X0Y225_ILOGIC_X0Y225_O = LIOB33_X0Y225_IOB_X0Y225_I;
  assign LIOI3_X0Y227_ILOGIC_X0Y228_O = LIOB33_X0Y227_IOB_X0Y228_I;
  assign LIOI3_X0Y227_ILOGIC_X0Y227_O = LIOB33_X0Y227_IOB_X0Y227_I;
  assign LIOI3_X0Y229_ILOGIC_X0Y230_O = LIOB33_X0Y229_IOB_X0Y230_I;
  assign LIOI3_X0Y229_ILOGIC_X0Y229_O = LIOB33_X0Y229_IOB_X0Y229_I;
  assign LIOI3_X0Y233_ILOGIC_X0Y234_O = LIOB33_X0Y233_IOB_X0Y234_I;
  assign LIOI3_X0Y235_ILOGIC_X0Y236_O = LIOB33_X0Y235_IOB_X0Y236_I;
  assign LIOI3_X0Y235_ILOGIC_X0Y235_O = LIOB33_X0Y235_IOB_X0Y235_I;
  assign LIOI3_X0Y239_ILOGIC_X0Y240_O = LIOB33_X0Y239_IOB_X0Y240_I;
  assign LIOI3_X0Y239_ILOGIC_X0Y239_O = LIOB33_X0Y239_IOB_X0Y239_I;
  assign LIOI3_X0Y241_ILOGIC_X0Y242_O = LIOB33_X0Y241_IOB_X0Y242_I;
  assign LIOI3_X0Y241_ILOGIC_X0Y241_O = LIOB33_X0Y241_IOB_X0Y241_I;
  assign LIOI3_SING_X0Y0_ILOGIC_X0Y0_O = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y99_ILOGIC_X0Y99_O = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_ILOGIC_X0Y149_O = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_O = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign LIOI3_SING_X0Y199_ILOGIC_X0Y199_O = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign LIOI3_SING_X0Y200_ILOGIC_X0Y200_O = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_O = LIOB33_X0Y19_IOB_X0Y20_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_O = LIOB33_X0Y19_IOB_X0Y19_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_O = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_O = LIOB33_X0Y81_IOB_X0Y81_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_O = LIOB33_X0Y93_IOB_X0Y94_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_O = LIOB33_X0Y93_IOB_X0Y93_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O = LIOB33_X0Y119_IOB_X0Y119_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O = LIOB33_X0Y131_IOB_X0Y132_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O = LIOB33_X0Y131_IOB_X0Y131_I;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_O = LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_D;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O = LIOB33_X0Y157_IOB_X0Y157_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_O = LIOB33_X0Y169_IOB_X0Y170_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_O = LIOB33_X0Y169_IOB_X0Y169_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_O = LIOB33_X0Y181_IOB_X0Y182_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_O = LIOB33_X0Y181_IOB_X0Y181_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_O = LIOB33_X0Y193_IOB_X0Y194_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_O = LIOB33_X0Y193_IOB_X0Y193_I;
  assign LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y208_O = LIOB33_X0Y207_IOB_X0Y208_I;
  assign LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y207_O = LIOB33_X0Y207_IOB_X0Y207_I;
  assign LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y220_O = LIOB33_X0Y219_IOB_X0Y220_I;
  assign LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y219_O = LIOB33_X0Y219_IOB_X0Y219_I;
  assign LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y232_O = LIOB33_X0Y231_IOB_X0Y232_I;
  assign LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y231_O = LIOB33_X0Y231_IOB_X0Y231_I;
  assign LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y243_O = LIOB33_X0Y243_IOB_X0Y243_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_O = LIOB33_X0Y13_IOB_X0Y14_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_O = LIOB33_X0Y13_IOB_X0Y13_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_O = LIOB33_X0Y87_IOB_X0Y88_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_O = LIOB33_X0Y87_IOB_X0Y87_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O = LIOB33_X0Y163_IOB_X0Y164_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_O = LIOB33_X0Y187_IOB_X0Y188_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_O = LIOB33_X0Y187_IOB_X0Y187_I;
  assign LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y214_O = LIOB33_X0Y213_IOB_X0Y214_I;
  assign LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y213_O = LIOB33_X0Y213_IOB_X0Y213_I;
  assign LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y238_O = LIOB33_X0Y237_IOB_X0Y238_I;
  assign LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y237_O = LIOB33_X0Y237_IOB_X0Y237_I;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_OQ = LIOB33_X0Y77_IOB_X0Y78_I;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_OQ = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_OQ = LIOB33_X0Y79_IOB_X0Y80_I;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_TQ = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_OQ = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_TQ = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_OQ = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_TQ = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_OQ = CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_OQ = LIOB33_X0Y83_IOB_X0Y84_I;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_TQ = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_OQ = LIOB33_X0Y83_IOB_X0Y83_I;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_TQ = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_OQ = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_TQ = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_OQ = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_OQ = LIOB33_X0Y89_IOB_X0Y90_I;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_OQ = LIOB33_X0Y87_IOB_X0Y88_I;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_OQ = LIOB33_X0Y91_IOB_X0Y92_I;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_OQ = LIOB33_X0Y91_IOB_X0Y91_I;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_OQ = CLBLL_L_X2Y189_SLICE_X0Y189_AO6;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_OQ = LIOB33_X0Y95_IOB_X0Y95_I;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_OQ = CLBLM_L_X44Y158_SLICE_X66Y158_BO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_OQ = LIOB33_X0Y95_IOB_X0Y96_I;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_OQ = LIOB33_X0Y97_IOB_X0Y97_I;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_OQ = CLBLM_L_X44Y152_SLICE_X66Y152_AO6;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_TQ = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_OQ = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_TQ = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_OQ = LIOB33_X0Y97_IOB_X0Y98_I;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_OQ = CLBLL_L_X2Y208_SLICE_X0Y208_AO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_OQ = LIOB33_X0Y109_IOB_X0Y109_I;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_OQ = CLBLL_L_X2Y187_SLICE_X0Y187_AO6;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_OQ = CLBLL_L_X2Y189_SLICE_X1Y189_AO6;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_OQ = CLBLL_L_X2Y194_SLICE_X0Y194_AO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_OQ = LIOB33_X0Y109_IOB_X0Y110_I;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_OQ = LIOB33_X0Y113_IOB_X0Y113_I;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_OQ = LIOB33_X0Y111_IOB_X0Y112_I;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_OQ = LIOB33_X0Y115_IOB_X0Y115_I;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_OQ = LIOB33_X0Y113_IOB_X0Y114_I;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_TQ = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_OQ = LIOB33_X0Y119_IOB_X0Y120_I;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_TQ = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_OQ = LIOB33_X0Y117_IOB_X0Y118_I;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_TQ = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_OQ = LIOB33_X0Y121_IOB_X0Y122_I;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_TQ = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_OQ = LIOB33_X0Y121_IOB_X0Y121_I;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_OQ = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_OQ = LIOB33_X0Y81_IOB_X0Y81_I;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_OQ = CLBLL_L_X2Y189_SLICE_X1Y189_AO6;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_OQ = LIOB33_X0Y203_IOB_X0Y204_I;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_OQ = LIOB33_X0Y203_IOB_X0Y203_I;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_OQ = CLBLL_L_X2Y192_SLICE_X0Y192_BO6;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_OQ = LIOB33_X0Y205_IOB_X0Y205_I;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_OQ = CLBLL_L_X2Y192_SLICE_X0Y192_CO6;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_OQ = CLBLL_L_X2Y193_SLICE_X0Y193_BO6;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_OQ = CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_OQ = CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_OQ = CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_OQ = CLBLL_L_X2Y154_SLICE_X0Y154_AO6;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_OQ = CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_OQ = CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_OQ = CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_OQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_TQ = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_OQ = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_TQ = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = CLBLM_R_X59Y133_SLICE_X88Y133_AO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_OQ = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_OQ = LIOB33_X0Y183_IOB_X0Y184_I;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_OQ = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_OQ = LIOB33_X0Y229_IOB_X0Y230_I;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_OQ = LIOB33_X0Y9_IOB_X0Y10_I;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_OQ = LIOB33_X0Y103_IOB_X0Y104_I;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_OQ = LIOB33_X0Y195_IOB_X0Y195_I;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_OQ = CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_OQ = CLBLL_L_X2Y149_SLICE_X0Y149_AO5;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_TQ = 1'b1;
  assign RIOI3_X105Y151_ILOGIC_X1Y152_O = RIOB33_X105Y151_IOB_X1Y152_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y151_O = RIOB33_X105Y151_IOB_X1Y151_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y154_O = RIOB33_X105Y153_IOB_X1Y154_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y153_O = RIOB33_X105Y153_IOB_X1Y153_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y156_O = RIOB33_X105Y155_IOB_X1Y156_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y155_O = RIOB33_X105Y155_IOB_X1Y155_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y159_O = RIOB33_X105Y159_IOB_X1Y159_I;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_R_X59Y159_SLICE_X88Y159_AO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X44Y158_SLICE_X66Y158_AO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X44Y158_SLICE_X66Y158_BO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = CLBLM_R_X47Y158_SLICE_X72Y158_AO5;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = LIOB33_X0Y19_IOB_X0Y19_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = LIOB33_X0Y21_IOB_X0Y21_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_X0Y19_IOB_X0Y20_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = LIOB33_X0Y25_IOB_X0Y25_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = LIOB33_X0Y23_IOB_X0Y24_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = LIOB33_X0Y27_IOB_X0Y28_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = LIOB33_X0Y27_IOB_X0Y27_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = LIOB33_X0Y53_IOB_X0Y53_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLL_L_X2Y193_SLICE_X0Y193_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_OQ = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ = 1'b1;
  assign RIOI3_SING_X105Y150_ILOGIC_X1Y150_O = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = LIOB33_X0Y241_IOB_X0Y242_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_OQ = LIOB33_X0Y81_IOB_X0Y82_I;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_OQ = CLBLL_L_X2Y210_SLICE_X0Y210_AO6;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ = LIOB33_X0Y93_IOB_X0Y94_I;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ = LIOB33_X0Y93_IOB_X0Y93_I;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ = CLBLL_L_X2Y193_SLICE_X0Y193_AO6;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ = CLBLL_L_X2Y210_SLICE_X0Y210_AO6;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_OQ = LIOB33_X0Y117_IOB_X0Y117_I;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_OQ = LIOB33_X0Y115_IOB_X0Y116_I;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ = LIOB33_X0Y201_IOB_X0Y202_I;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ = LIOB33_X0Y201_IOB_X0Y201_I;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ = CLBLM_R_X67Y130_SLICE_X100Y130_AO6;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = CLBLM_R_X59Y133_SLICE_X88Y133_AO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ = LIOB33_X0Y1_IOB_X0Y1_I;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ = LIOB33_X0Y217_IOB_X0Y217_I;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_O = RIOB33_X105Y157_IOB_X1Y158_I;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_O = RIOB33_X105Y157_IOB_X1Y157_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = LIOB33_X0Y23_IOB_X0Y23_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = LIOB33_X0Y21_IOB_X0Y22_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X44Y152_SLICE_X66Y152_AO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ = LIOB33_X0Y87_IOB_X0Y87_I;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ = LIOB33_X0Y85_IOB_X0Y86_I;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ = LIOB33_X0Y111_IOB_X0Y111_I;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ = CLBLL_L_X2Y192_SLICE_X0Y192_AO6;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ = CLBLL_L_X2Y193_SLICE_X0Y193_BO6;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ = CLBLL_L_X2Y192_SLICE_X0Y192_BO6;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ = LIOB33_X0Y135_IOB_X0Y135_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ = LIOB33_X0Y135_IOB_X0Y135_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_R_X47Y158_SLICE_X72Y158_AO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X44Y158_SLICE_X66Y158_AO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y176_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign RIOB33_X105Y175_IOB_X1Y175_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOB33_SING_X105Y149_IOB_X1Y149_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_D = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = LIOB33_X0Y25_IOB_X0Y25_I;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_D1 = LIOB33_X0Y183_IOB_X0Y184_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_D1 = LIOB33_X0Y203_IOB_X0Y204_I;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_T1 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_D1 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = LIOB33_X0Y23_IOB_X0Y24_I;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_A1 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_A2 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_A3 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_A4 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_A5 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_A6 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_T1 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_D1 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_T1 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_B1 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_B2 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_B3 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_B4 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_B5 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_B6 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_D1 = LIOB33_X0Y203_IOB_X0Y203_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_T1 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_C1 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_C2 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_C3 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_C4 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_C5 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_C6 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_D1 = LIOB33_X0Y97_IOB_X0Y98_I;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_T1 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_D1 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_D2 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_D3 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_D4 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A1 = LIOB33_X0Y209_IOB_X0Y209_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A2 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A3 = LIOB33_X0Y207_IOB_X0Y208_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A4 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A5 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A6 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X67Y158_D6 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_A1 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B6 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_A2 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_A3 = LIOB33_X0Y217_IOB_X0Y218_I;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_A5 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C6 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_B2 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_B3 = LIOB33_X0Y217_IOB_X0Y218_I;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_B4 = CLBLM_R_X47Y158_SLICE_X72Y158_BO6;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_B5 = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_B6 = 1'b1;
  assign RIOB33_X105Y57_IOB_X1Y58_O = LIOB33_X0Y81_IOB_X0Y82_I;
  assign RIOB33_X105Y57_IOB_X1Y57_O = CLBLL_L_X2Y210_SLICE_X0Y210_AO6;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D6 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_C3 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_C4 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_D1 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_D2 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_D3 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_D4 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_D5 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_D6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A6 = 1'b1;
  assign RIOB33_X105Y117_IOB_X1Y117_O = CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  assign RIOB33_X105Y117_IOB_X1Y118_O = CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C6 = 1'b1;
  assign LIOI3_X0Y217_ILOGIC_X0Y218_D = LIOB33_X0Y217_IOB_X0Y218_I;
  assign LIOI3_X0Y217_ILOGIC_X0Y217_D = LIOB33_X0Y217_IOB_X0Y217_I;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D6 = 1'b1;
  assign LIOI3_X0Y185_ILOGIC_X0Y186_D = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y185_D = LIOB33_X0Y185_IOB_X0Y185_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_D = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_D = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOB33_X105Y177_IOB_X1Y178_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign RIOB33_X105Y177_IOB_X1Y177_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = LIOB33_X0Y241_IOB_X0Y242_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y96_D = LIOB33_X0Y95_IOB_X0Y96_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y95_D = LIOB33_X0Y95_IOB_X0Y95_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y4_D = LIOB33_X0Y3_IOB_X0Y4_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y3_D = LIOB33_X0Y3_IOB_X0Y3_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_D = LIOB33_X0Y13_IOB_X0Y14_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_D = LIOB33_X0Y13_IOB_X0Y13_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_A1 = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_A2 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_A3 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_A4 = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_A5 = LIOB33_X0Y167_IOB_X0Y168_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_A6 = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_B1 = LIOB33_X0Y15_IOB_X0Y15_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_B2 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_B3 = CLBLL_L_X2Y170_SLICE_X0Y170_AO6;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_B4 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_B5 = CLBLL_L_X2Y165_SLICE_X0Y165_AO6;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_B6 = CLBLL_L_X2Y165_SLICE_X0Y165_CO6;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_C1 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_C2 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_C3 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_C4 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_C5 = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_C6 = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_D1 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_D2 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_D3 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_D4 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_D5 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X0Y165_D6 = 1'b1;
  assign LIOI3_SING_X0Y199_ILOGIC_X0Y199_D = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_A1 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_A2 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_A3 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_A4 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_A5 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_B1 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_B2 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_B3 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_B4 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_B5 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_B6 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_C1 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_C2 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_C3 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_C4 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_C5 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_C6 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_D1 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_D2 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_D3 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_D4 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_D5 = 1'b1;
  assign CLBLL_L_X2Y165_SLICE_X1Y165_D6 = 1'b1;
  assign RIOB33_X105Y59_IOB_X1Y60_O = LIOB33_X0Y83_IOB_X0Y84_I;
  assign RIOB33_X105Y59_IOB_X1Y59_O = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_A1 = LIOB33_X0Y219_IOB_X0Y219_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_A2 = LIOB33_X0Y231_IOB_X0Y231_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_A3 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_A4 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_A5 = LIOB33_X0Y197_IOB_X0Y197_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_A6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign RIOB33_X105Y119_IOB_X1Y119_O = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign RIOB33_X105Y119_IOB_X1Y120_O = CLBLM_R_X67Y130_SLICE_X100Y130_AO6;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_B1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_B2 = LIOB33_X0Y237_IOB_X0Y238_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_B3 = LIOB33_X0Y191_IOB_X0Y192_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_B4 = LIOB33_X0Y225_IOB_X0Y226_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_B5 = LIOB33_X0Y213_IOB_X0Y214_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_B6 = CLBLL_L_X2Y210_SLICE_X0Y210_BO6;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_C1 = LIOB33_X0Y191_IOB_X0Y192_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_C2 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_C3 = LIOB33_X0Y213_IOB_X0Y214_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_C4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_C5 = LIOB33_X0Y237_IOB_X0Y238_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_C6 = LIOB33_X0Y225_IOB_X0Y226_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_D1 = LIOB33_X0Y231_IOB_X0Y231_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_D2 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_D3 = LIOB33_X0Y197_IOB_X0Y197_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_D4 = CLBLL_L_X2Y187_SLICE_X0Y187_AO5;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_D5 = LIOB33_X0Y219_IOB_X0Y219_I;
  assign CLBLL_L_X2Y192_SLICE_X0Y192_D6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign RIOB33_X105Y179_IOB_X1Y180_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOB33_X105Y179_IOB_X1Y179_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_A1 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_A2 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_A3 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_A4 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_A5 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_A6 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_B1 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_B2 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_B3 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_B4 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_B5 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_B6 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_C1 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_C2 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_C3 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_C4 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_C5 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_C6 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_D1 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_D2 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_D3 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_D4 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_D5 = 1'b1;
  assign CLBLL_L_X2Y192_SLICE_X1Y192_D6 = 1'b1;
  assign LIOI3_SING_X0Y200_ILOGIC_X0Y200_D = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign RIOB33_X105Y61_IOB_X1Y62_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOB33_X105Y61_IOB_X1Y61_O = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOB33_X105Y121_IOB_X1Y122_O = CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  assign RIOB33_X105Y121_IOB_X1Y121_O = CLBLL_L_X2Y154_SLICE_X0Y154_AO6;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_A1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_A2 = LIOB33_X0Y211_IOB_X0Y211_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_A3 = LIOB33_X0Y189_IOB_X0Y190_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_A4 = LIOB33_X0Y223_IOB_X0Y223_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_A5 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_A6 = LIOB33_X0Y235_IOB_X0Y235_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_B1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_B2 = CLBLL_L_X2Y208_SLICE_X0Y208_BO6;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_B3 = LIOB33_X0Y211_IOB_X0Y211_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_B4 = LIOB33_X0Y223_IOB_X0Y223_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_B5 = LIOB33_X0Y189_IOB_X0Y190_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_B6 = LIOB33_X0Y235_IOB_X0Y235_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = LIOB33_X0Y27_IOB_X0Y28_I;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_D1 = LIOB33_X0Y229_IOB_X0Y230_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_C1 = LIOB33_X0Y191_IOB_X0Y192_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_C2 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_C3 = LIOB33_X0Y213_IOB_X0Y214_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_C4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_C5 = LIOB33_X0Y237_IOB_X0Y238_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_C6 = LIOB33_X0Y225_IOB_X0Y226_I;
  assign RIOB33_X105Y181_IOB_X1Y181_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOB33_X105Y181_IOB_X1Y182_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_D1 = CLBLL_L_X2Y192_SLICE_X0Y192_BO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_T1 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_D1 = LIOB33_X0Y189_IOB_X0Y190_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_D2 = LIOB33_X0Y227_IOB_X0Y227_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_D3 = LIOB33_X0Y223_IOB_X0Y223_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_D4 = CLBLL_L_X2Y187_SLICE_X0Y187_AO5;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_D5 = LIOB33_X0Y211_IOB_X0Y211_I;
  assign CLBLL_L_X2Y193_SLICE_X0Y193_D6 = LIOB33_X0Y235_IOB_X0Y235_I;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_D1 = CLBLL_L_X2Y208_SLICE_X0Y208_AO6;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_D1 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_D1 = LIOB33_X0Y9_IOB_X0Y10_I;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_D1 = LIOB33_X0Y205_IOB_X0Y205_I;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_T1 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_D1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_R_X47Y158_SLICE_X72Y158_AO5;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_T1 = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_A1 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_A2 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_A3 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_A4 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_A5 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_A6 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_D1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_B1 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_B2 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_B3 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_B4 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_B5 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X44Y158_SLICE_X66Y158_AO6;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_C1 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_C2 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_C3 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_C4 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_C5 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X44Y152_SLICE_X66Y152_AO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_D1 = CLBLL_L_X2Y210_SLICE_X0Y210_AO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_D1 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_D2 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_D3 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_D4 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_D5 = 1'b1;
  assign CLBLL_L_X2Y193_SLICE_X1Y193_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_T1 = 1'b1;
  assign LIOI3_X0Y221_ILOGIC_X0Y222_D = LIOB33_X0Y221_IOB_X0Y222_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y190_D = LIOB33_X0Y189_IOB_X0Y190_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y189_D = LIOB33_X0Y189_IOB_X0Y189_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_D = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_D = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y98_D = LIOB33_X0Y97_IOB_X0Y98_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y97_D = LIOB33_X0Y97_IOB_X0Y97_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign RIOB33_X105Y63_IOB_X1Y64_O = LIOB33_X0Y87_IOB_X0Y87_I;
  assign RIOB33_X105Y63_IOB_X1Y63_O = LIOB33_X0Y85_IOB_X0Y86_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_D = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_D = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D = LIOB33_X0Y131_IOB_X0Y132_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D = LIOB33_X0Y131_IOB_X0Y131_I;
  assign RIOB33_X105Y123_IOB_X1Y124_O = CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  assign RIOB33_X105Y123_IOB_X1Y123_O = CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  assign RIOB33_X105Y183_IOB_X1Y184_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_A1 = 1'b1;
  assign RIOB33_X105Y183_IOB_X1Y183_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_A2 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_A3 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_A1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_A2 = LIOB33_X0Y219_IOB_X0Y220_I;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_A3 = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_A4 = LIOB33_X0Y197_IOB_X0Y198_I;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_A5 = LIOB33_X0Y231_IOB_X0Y232_I;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_A6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_B1 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_B2 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_B3 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_B1 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_B2 = LIOB33_X0Y219_IOB_X0Y220_I;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_B3 = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_B4 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_B5 = LIOB33_X0Y231_IOB_X0Y232_I;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_B6 = LIOB33_X0Y197_IOB_X0Y198_I;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_B4 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_B6 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_C3 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_C1 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_C2 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_C3 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_C4 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_C5 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_C6 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_C4 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_C5 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_C6 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_D1 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_D2 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_D3 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_D4 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_D1 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_D2 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_D3 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_D4 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_D5 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X0Y194_D6 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_D5 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_D6 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_A1 = LIOB33_X0Y217_IOB_X0Y217_I;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_A2 = LIOB33_X0Y1_IOB_X0Y1_I;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_A4 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_A5 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_A6 = LIOB33_X0Y195_IOB_X0Y195_I;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_B1 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_B2 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_B3 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_B4 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_B5 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_B6 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_C1 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_C2 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_C3 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_C4 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_C5 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_A1 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_A2 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_A3 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_A4 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_A5 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_A6 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_C6 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_B1 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_B2 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_B3 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_B4 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_B5 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_B6 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_D1 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_D2 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_D3 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_C1 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_C2 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_C3 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_C4 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_C5 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_C6 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_D1 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_D2 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_D3 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_D4 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_D5 = 1'b1;
  assign CLBLL_L_X2Y194_SLICE_X1Y194_D6 = 1'b1;
  assign RIOB33_X105Y65_IOB_X1Y66_O = LIOB33_X0Y89_IOB_X0Y90_I;
  assign RIOB33_X105Y65_IOB_X1Y65_O = LIOB33_X0Y87_IOB_X0Y88_I;
  assign RIOB33_X105Y125_IOB_X1Y126_O = CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  assign RIOB33_X105Y125_IOB_X1Y125_O = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_A1 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_A2 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_A3 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_A4 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_A5 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_A6 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_B1 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_B2 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_B3 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_B4 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_B5 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_B6 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_C1 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_C2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A1 = CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A2 = LIOB33_X0Y195_IOB_X0Y196_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A3 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A4 = LIOB33_X0Y187_IOB_X0Y188_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A5 = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A6 = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_C3 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_C4 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_C5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_D1 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_D2 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_D3 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_D4 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_D5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B3 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B4 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B5 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C1 = CLBLL_L_X2Y142_SLICE_X0Y142_AO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C2 = CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C3 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C5 = CLBLL_L_X2Y142_SLICE_X0Y142_DO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C6 = CLBLL_L_X2Y142_SLICE_X0Y142_BO6;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_A1 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_A2 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_A5 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_A3 = CLBLL_L_X2Y165_SLICE_X0Y165_BO6;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_A4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D1 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D2 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D3 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D4 = LIOB33_X0Y207_IOB_X0Y207_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_B1 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_B2 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_B3 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_B4 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_B5 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_B6 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_C1 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_C2 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_C3 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_C4 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_C5 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_C6 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_D1 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_D2 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_D3 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_D4 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_D5 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_D6 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A6 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B6 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C6 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D6 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_D1 = CLBLL_L_X2Y192_SLICE_X0Y192_CO6;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_T1 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_D1 = CLBLL_L_X2Y187_SLICE_X0Y187_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_T1 = 1'b1;
  assign RIOB33_X105Y67_IOB_X1Y68_O = LIOB33_X0Y91_IOB_X0Y92_I;
  assign RIOB33_X105Y67_IOB_X1Y67_O = LIOB33_X0Y91_IOB_X0Y91_I;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_D1 = LIOB33_X0Y195_IOB_X0Y195_I;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_D1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_D1 = CLBLL_L_X2Y193_SLICE_X0Y193_BO6;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_T1 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_T1 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_D1 = CLBLL_L_X2Y189_SLICE_X1Y189_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_T1 = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1 = LIOB33_X0Y93_IOB_X0Y94_I;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign RIOB33_X105Y127_IOB_X1Y128_O = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign RIOB33_X105Y127_IOB_X1Y127_O = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y188_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOB33_X105Y187_IOB_X1Y187_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y223_ILOGIC_X0Y224_D = LIOB33_X0Y223_IOB_X0Y224_I;
  assign LIOI3_X0Y223_ILOGIC_X0Y223_D = LIOB33_X0Y223_IOB_X0Y223_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y192_D = LIOB33_X0Y191_IOB_X0Y192_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y191_D = LIOB33_X0Y191_IOB_X0Y191_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_D = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_D = LIOB33_X0Y161_IOB_X0Y161_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_D = LIOB33_X0Y129_IOB_X0Y130_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_D = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_D = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_D = LIOB33_X0Y27_IOB_X0Y27_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_D = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D = LIOB33_X0Y7_IOB_X0Y7_I;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_A1 = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_A2 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_A3 = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_A4 = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_A5 = LIOB33_X0Y169_IOB_X0Y170_I;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_A6 = 1'b1;
  assign RIOB33_X105Y69_IOB_X1Y70_O = LIOB33_X0Y93_IOB_X0Y94_I;
  assign RIOB33_X105Y69_IOB_X1Y69_O = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_B1 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_B2 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_B3 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_B4 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_B5 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_B6 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_C1 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_C2 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_C3 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_C4 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_C5 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_C6 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_D1 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_D2 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_D3 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_D4 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_D5 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X0Y170_D6 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_A4 = LIOB33_X0Y165_IOB_X0Y165_I;
  assign RIOB33_X105Y129_IOB_X1Y130_O = CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  assign RIOB33_X105Y129_IOB_X1Y129_O = CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_A6 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_A1 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_A2 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_A3 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_A4 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_A5 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_A6 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_B1 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_B2 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_B3 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_B4 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_B5 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_B6 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_B1 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_C1 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_C2 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_C3 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_C4 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_C5 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_C6 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y190_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign RIOB33_X105Y189_IOB_X1Y189_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_D1 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_D2 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_D3 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_D4 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_D5 = 1'b1;
  assign CLBLL_L_X2Y170_SLICE_X1Y170_D6 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_C2 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_C5 = 1'b1;
  assign CLBLM_L_X44Y158_SLICE_X66Y158_C6 = 1'b1;
  assign RIOB33_X105Y71_IOB_X1Y72_O = CLBLL_L_X2Y189_SLICE_X0Y189_AO6;
  assign RIOB33_X105Y71_IOB_X1Y71_O = LIOB33_X0Y95_IOB_X0Y95_I;
  assign RIOB33_X105Y131_IOB_X1Y132_O = CLBLM_R_X59Y133_SLICE_X88Y133_AO6;
  assign RIOB33_X105Y131_IOB_X1Y131_O = 1'b0;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOB33_X105Y191_IOB_X1Y191_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A1 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A2 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A4 = CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A5 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A6 = CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_D1 = CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B1 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_D1 = CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B2 = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B4 = LIOB33_X0Y205_IOB_X0Y206_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B5 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_T1 = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_D1 = CLBLL_L_X2Y194_SLICE_X0Y194_AO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C2 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C3 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_T1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C6 = LIOB33_X0Y205_IOB_X0Y206_I;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_D1 = CLBLL_L_X2Y149_SLICE_X0Y149_AO5;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_D1 = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D1 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D2 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D3 = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D4 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D6 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_D1 = CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_T1 = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_T1 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_T1 = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_D1 = CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1 = CLBLL_L_X2Y193_SLICE_X0Y193_AO6;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1 = CLBLL_L_X2Y210_SLICE_X0Y210_AO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D6 = 1'b1;
  assign RIOB33_X105Y73_IOB_X1Y74_O = CLBLM_L_X44Y158_SLICE_X66Y158_BO6;
  assign RIOB33_X105Y73_IOB_X1Y73_O = LIOB33_X0Y95_IOB_X0Y96_I;
  assign LIOI3_X0Y225_ILOGIC_X0Y226_D = LIOB33_X0Y225_IOB_X0Y226_I;
  assign LIOI3_X0Y225_ILOGIC_X0Y225_D = LIOB33_X0Y225_IOB_X0Y225_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y196_D = LIOB33_X0Y195_IOB_X0Y196_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y195_D = LIOB33_X0Y195_IOB_X0Y195_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_D = LIOB33_X0Y165_IOB_X0Y166_I;
  assign RIOB33_X105Y133_IOB_X1Y134_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOB33_X105Y133_IOB_X1Y133_O = CLBLM_R_X59Y133_SLICE_X88Y133_AO6;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_D = LIOB33_X0Y165_IOB_X0Y165_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_D = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_D = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_D = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_D = LIOB33_X0Y11_IOB_X0Y11_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X44Y152_SLICE_X66Y152_AO5;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_D = LIOB33_X0Y87_IOB_X0Y88_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_D = LIOB33_X0Y87_IOB_X0Y87_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D = LIOB33_X0Y157_IOB_X0Y157_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_D = LIOB33_X0Y19_IOB_X0Y20_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_D = LIOB33_X0Y19_IOB_X0Y19_I;
  assign RIOB33_X105Y75_IOB_X1Y76_O = LIOB33_X0Y97_IOB_X0Y97_I;
  assign RIOB33_X105Y75_IOB_X1Y75_O = CLBLM_L_X44Y152_SLICE_X66Y152_AO6;
  assign RIOB33_X105Y135_IOB_X1Y136_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOB33_X105Y135_IOB_X1Y135_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLL_L_X2Y193_SLICE_X0Y193_AO6;
  assign RIOB33_X105Y195_IOB_X1Y195_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A1 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A2 = CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A3 = CLBLL_L_X2Y134_SLICE_X0Y134_CO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A4 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A5 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A6 = LIOB33_X0Y205_IOB_X0Y206_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B3 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B5 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B6 = LIOB33_X0Y25_IOB_X0Y26_I;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C6 = 1'b1;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B1 = 1'b1;
  assign RIOB33_X105Y77_IOB_X1Y78_O = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign RIOB33_X105Y77_IOB_X1Y77_O = LIOB33_X0Y97_IOB_X0Y98_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D6 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOB33_X105Y137_IOB_X1Y138_O = LIOB33_X0Y135_IOB_X0Y135_I;
  assign RIOB33_X105Y137_IOB_X1Y137_O = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_B2 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_D1 = CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_T1 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_D1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_D1 = CLBLL_L_X2Y154_SLICE_X0Y154_AO6;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_T1 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign RIOB33_X105Y197_IOB_X1Y198_O = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOB33_X105Y197_IOB_X1Y197_O = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_T1 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_D1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_T1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_B3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_B4 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_T1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_B5 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_T1 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_T1 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_D4 = 1'b1;
  assign LIOI3_X0Y227_ILOGIC_X0Y228_D = LIOB33_X0Y227_IOB_X0Y228_I;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_D5 = 1'b1;
  assign LIOI3_X0Y227_ILOGIC_X0Y227_D = LIOB33_X0Y227_IOB_X0Y227_I;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_D6 = 1'b1;
  assign LIOI3_X0Y197_ILOGIC_X0Y198_D = LIOB33_X0Y197_IOB_X0Y198_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y197_D = LIOB33_X0Y197_IOB_X0Y197_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y168_D = LIOB33_X0Y167_IOB_X0Y168_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y136_D = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A1 = CLBLL_L_X2Y149_SLICE_X1Y149_AO5;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A2 = CLBLL_L_X2Y189_SLICE_X0Y189_CO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A3 = LIOB33_X0Y227_IOB_X0Y227_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A5 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A6 = CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_D = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B1 = CLBLL_L_X2Y149_SLICE_X1Y149_AO5;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B2 = CLBLL_L_X2Y192_SLICE_X0Y192_DO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B3 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B5 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B6 = CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C1 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C2 = LIOB33_X0Y205_IOB_X0Y206_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C3 = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C4 = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C5 = CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C6 = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign RIOI3_X105Y151_ILOGIC_X1Y152_D = RIOB33_X105Y151_IOB_X1Y152_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y151_D = RIOB33_X105Y151_IOB_X1Y151_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_D = LIOB33_X0Y15_IOB_X0Y16_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_D = LIOB33_X0Y15_IOB_X0Y15_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D1 = CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D3 = CLBLL_L_X2Y149_SLICE_X0Y149_BO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D4 = CLBLL_L_X2Y149_SLICE_X0Y149_CO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D5 = CLBLL_L_X2Y149_SLICE_X0Y149_DO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D6 = CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_D = LIOB33_X0Y169_IOB_X0Y170_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_D = LIOB33_X0Y169_IOB_X0Y169_I;
  assign RIOB33_X105Y79_IOB_X1Y80_O = CLBLL_L_X2Y208_SLICE_X0Y208_AO6;
  assign RIOB33_X105Y79_IOB_X1Y79_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_D1 = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A6 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_A4 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_A5 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_A5 = CLBLL_L_X2Y154_SLICE_X0Y154_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B6 = 1'b1;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_T1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C6 = 1'b1;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_D = LIOB33_X0Y145_IOB_X0Y146_I;
  assign RIOB33_X105Y139_IOB_X1Y140_O = LIOB33_X0Y183_IOB_X0Y184_I;
  assign RIOB33_X105Y139_IOB_X1Y139_O = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D6 = 1'b1;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_D = LIOB33_X0Y145_IOB_X0Y145_I;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1 = LIOB33_X0Y1_IOB_X0Y1_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A1 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A2 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A3 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A4 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A5 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A6 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B1 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B2 = CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B3 = CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B4 = CLBLL_L_X2Y193_SLICE_X0Y193_DO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B5 = CLBLL_L_X2Y210_SLICE_X0Y210_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B6 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_D = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C1 = CLBLL_L_X2Y149_SLICE_X0Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C2 = CLBLL_L_X2Y149_SLICE_X1Y149_CO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C3 = CLBLL_L_X2Y150_SLICE_X0Y150_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C4 = CLBLL_L_X2Y210_SLICE_X0Y210_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C5 = CLBLL_L_X2Y208_SLICE_X0Y208_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C6 = CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  assign RIOB33_X105Y81_IOB_X1Y82_O = CLBLL_L_X2Y193_SLICE_X0Y193_AO6;
  assign RIOB33_X105Y81_IOB_X1Y81_O = CLBLL_L_X2Y210_SLICE_X0Y210_AO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D1 = CLBLL_L_X2Y193_SLICE_X0Y193_AO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D2 = CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D3 = CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D5 = LIOB33_X0Y227_IOB_X0Y227_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D6 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = LIOB33_X0Y27_IOB_X0Y27_I;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1 = LIOB33_X0Y87_IOB_X0Y87_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A1 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A2 = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A3 = 1'b1;
  assign RIOB33_X105Y141_IOB_X1Y142_O = LIOB33_X0Y229_IOB_X0Y230_I;
  assign RIOB33_X105Y141_IOB_X1Y141_O = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A4 = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A5 = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A6 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B1 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B2 = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B3 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B4 = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B5 = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B6 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C1 = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C2 = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C3 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C4 = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C5 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C6 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_C1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_C2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D6 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_C3 = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_C6 = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1 = 1'b1;
  assign LIOI3_X0Y205_ILOGIC_X0Y206_D = LIOB33_X0Y205_IOB_X0Y206_I;
  assign LIOI3_X0Y205_ILOGIC_X0Y205_D = LIOB33_X0Y205_IOB_X0Y205_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_D1 = CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y185_IOB_X1Y186_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_T1 = 1'b1;
  assign RIOB33_X105Y185_IOB_X1Y185_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_D1 = CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_T1 = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_T1 = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_D1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1 = LIOB33_X0Y201_IOB_X0Y202_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A1 = CLBLL_L_X2Y193_SLICE_X0Y193_CO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A2 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A4 = CLBLL_L_X2Y189_SLICE_X0Y189_BO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A5 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A6 = CLBLL_L_X2Y189_SLICE_X0Y189_CO6;
  assign RIOB33_X105Y83_IOB_X1Y83_O = CLBLL_L_X2Y189_SLICE_X1Y189_AO6;
  assign RIOB33_X105Y83_IOB_X1Y84_O = CLBLL_L_X2Y187_SLICE_X0Y187_AO6;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B1 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B2 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B3 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B4 = CLBLL_L_X2Y189_SLICE_X0Y189_BO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B5 = LIOB33_X0Y205_IOB_X0Y206_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B6 = CLBLL_L_X2Y193_SLICE_X0Y193_CO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C2 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C3 = CLBLL_L_X2Y193_SLICE_X0Y193_CO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C6 = CLBLL_L_X2Y189_SLICE_X0Y189_BO6;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1 = LIOB33_X0Y201_IOB_X0Y201_I;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D6 = 1'b1;
  assign RIOB33_X105Y143_IOB_X1Y144_O = LIOB33_X0Y1_IOB_X0Y1_I;
  assign RIOB33_X105Y143_IOB_X1Y143_O = LIOB33_X0Y217_IOB_X0Y217_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A6 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B6 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C6 = 1'b1;
  assign LIOI3_X0Y229_ILOGIC_X0Y230_D = LIOB33_X0Y229_IOB_X0Y230_I;
  assign LIOI3_X0Y229_ILOGIC_X0Y229_D = LIOB33_X0Y229_IOB_X0Y229_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D1 = 1'b1;
  assign LIOI3_X0Y201_ILOGIC_X0Y202_D = LIOB33_X0Y201_IOB_X0Y202_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D4 = 1'b1;
  assign LIOI3_X0Y201_ILOGIC_X0Y201_D = LIOB33_X0Y201_IOB_X0Y201_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D6 = 1'b1;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_D = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y140_D = LIOB33_X0Y139_IOB_X0Y140_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y139_D = LIOB33_X0Y139_IOB_X0Y139_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y154_D = RIOB33_X105Y153_IOB_X1Y154_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y153_D = RIOB33_X105Y153_IOB_X1Y153_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_D = LIOB33_X0Y17_IOB_X0Y18_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_D = LIOB33_X0Y17_IOB_X0Y17_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_D = LIOB33_X0Y181_IOB_X0Y182_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_D = LIOB33_X0Y181_IOB_X0Y181_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1 = 1'b1;
  assign RIOB33_X105Y85_IOB_X1Y86_O = CLBLL_L_X2Y194_SLICE_X0Y194_AO6;
  assign RIOB33_X105Y85_IOB_X1Y85_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A1 = CLBLL_L_X2Y193_SLICE_X0Y193_CO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A2 = CLBLL_L_X2Y193_SLICE_X0Y193_AO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A3 = CLBLL_L_X2Y208_SLICE_X0Y208_BO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A4 = CLBLL_L_X2Y189_SLICE_X0Y189_BO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A5 = CLBLL_L_X2Y210_SLICE_X0Y210_BO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A6 = CLBLL_L_X2Y210_SLICE_X0Y210_CO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B1 = CLBLL_L_X2Y193_SLICE_X0Y193_CO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B2 = CLBLL_L_X2Y187_SLICE_X0Y187_BO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B3 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B4 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B6 = CLBLL_L_X2Y210_SLICE_X0Y210_CO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C1 = CLBLL_L_X2Y151_SLICE_X0Y151_AO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C3 = LIOB33_X0Y179_IOB_X0Y180_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C5 = CLBLL_L_X2Y187_SLICE_X0Y187_BO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C6 = 1'b1;
  assign RIOB33_X105Y145_IOB_X1Y146_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign RIOB33_X105Y145_IOB_X1Y145_O = LIOB33_X0Y195_IOB_X0Y195_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D1 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D6 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A1 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A6 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B1 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B6 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C1 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C6 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D1 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D6 = 1'b1;
  assign RIOB33_X105Y87_IOB_X1Y88_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign RIOB33_X105Y87_IOB_X1Y87_O = CLBLL_L_X2Y192_SLICE_X0Y192_AO6;
  assign RIOB33_X105Y147_IOB_X1Y148_O = CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  assign RIOB33_X105Y147_IOB_X1Y147_O = CLBLL_L_X2Y149_SLICE_X0Y149_AO5;
  assign RIOI3_SING_X105Y150_ILOGIC_X1Y150_D = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_D1 = CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_D1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_T1 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_D1 = LIOB33_X0Y89_IOB_X0Y90_I;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_D1 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_T1 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_D1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_T1 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_D1 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1 = CLBLM_R_X67Y130_SLICE_X100Y130_AO6;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1 = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1 = 1'b1;
  assign LIOI3_X0Y233_ILOGIC_X0Y234_D = LIOB33_X0Y233_IOB_X0Y234_I;
  assign LIOI3_X0Y203_ILOGIC_X0Y204_D = LIOB33_X0Y203_IOB_X0Y204_I;
  assign LIOI3_X0Y203_ILOGIC_X0Y203_D = LIOB33_X0Y203_IOB_X0Y203_I;
  assign RIOB33_X105Y89_IOB_X1Y90_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign RIOB33_X105Y89_IOB_X1Y89_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_D = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_D = LIOB33_X0Y173_IOB_X0Y173_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_D = LIOB33_X0Y141_IOB_X0Y142_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_D = LIOB33_X0Y141_IOB_X0Y141_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y80_D = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y156_D = RIOB33_X105Y155_IOB_X1Y156_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y155_D = RIOB33_X105Y155_IOB_X1Y155_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = LIOB33_X0Y241_IOB_X0Y242_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_D = LIOB33_X0Y21_IOB_X0Y22_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_D = LIOB33_X0Y21_IOB_X0Y21_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D = LIOB33_X0Y163_IOB_X0Y164_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_D = LIOB33_X0Y193_IOB_X0Y194_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_D = LIOB33_X0Y193_IOB_X0Y193_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign RIOB33_X105Y91_IOB_X1Y92_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign RIOB33_X105Y91_IOB_X1Y91_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A1 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A3 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A4 = CLBLL_L_X2Y154_SLICE_X0Y154_BO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A5 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A6 = LIOB33_X0Y177_IOB_X0Y178_I;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B1 = LIOB33_X0Y207_IOB_X0Y208_I;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B2 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B3 = LIOB33_X0Y209_IOB_X0Y209_I;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B5 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B6 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C6 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D6 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A6 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B6 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C6 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D6 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_A1 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_A2 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_A3 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_A4 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_A5 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_A6 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_B1 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_B2 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_B3 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_B4 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_B5 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_B6 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_C1 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_C2 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_C3 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_C4 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_C5 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_C6 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_A5 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_A6 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_D1 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_D2 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_D3 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_D4 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_D5 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X73Y158_D6 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_A1 = LIOB33_X0Y229_IOB_X0Y230_I;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_A2 = LIOB33_X0Y241_IOB_X0Y242_I;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_A3 = CLBLM_R_X47Y145_SLICE_X72Y145_AO6;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_A4 = LIOB33_X0Y183_IOB_X0Y184_I;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_A5 = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_A6 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_B1 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_B2 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_B3 = CLBLM_R_X47Y145_SLICE_X72Y145_AO6;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_B4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_B5 = CLBLM_R_X47Y158_SLICE_X72Y158_AO6;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_B6 = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_C1 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_C2 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_C3 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_C4 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_C5 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_C6 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_B5 = 1'b1;
  assign RIOB33_X105Y93_IOB_X1Y94_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign RIOB33_X105Y93_IOB_X1Y93_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_R_X59Y159_SLICE_X88Y159_AO6;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_D1 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_D2 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_D3 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_D4 = 1'b1;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_D5 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_D1 = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign CLBLM_R_X47Y158_SLICE_X72Y158_D6 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_D1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_C1 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_T1 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_C2 = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_D1 = LIOB33_X0Y91_IOB_X0Y92_I;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_T1 = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_D1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_D1 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = CLBLM_R_X59Y133_SLICE_X88Y133_AO6;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A2 = LIOB33_X0Y13_IOB_X0Y14_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A5 = RIOB33_X105Y155_IOB_X1Y156_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A6 = LIOB33_X0Y5_IOB_X0Y5_I;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = 1'b0;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B6 = 1'b1;
  assign LIOI3_X0Y235_ILOGIC_X0Y235_D = LIOB33_X0Y235_IOB_X0Y235_I;
  assign LIOI3_X0Y235_ILOGIC_X0Y236_D = LIOB33_X0Y235_IOB_X0Y236_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C6 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_A1 = LIOB33_X0Y213_IOB_X0Y213_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_A2 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_A3 = LIOB33_X0Y225_IOB_X0Y225_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_A4 = LIOB33_X0Y237_IOB_X0Y237_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_A5 = LIOB33_X0Y191_IOB_X0Y191_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_A6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_B3 = LIOB33_X0Y191_IOB_X0Y191_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_B4 = LIOB33_X0Y237_IOB_X0Y237_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_B5 = LIOB33_X0Y225_IOB_X0Y225_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_B6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_B1 = LIOB33_X0Y213_IOB_X0Y213_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D5 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D6 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_C1 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_C2 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_C3 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_C4 = 1'b1;
  assign LIOI3_X0Y83_ILOGIC_X0Y84_D = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_C5 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_C6 = 1'b1;
  assign LIOI3_X0Y83_ILOGIC_X0Y83_D = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_D1 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_D2 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_D3 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_D4 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_D5 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X0Y208_D6 = 1'b1;
  assign RIOI3_X105Y159_ILOGIC_X1Y159_D = RIOB33_X105Y159_IOB_X1Y159_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_D = LIOB33_X0Y23_IOB_X0Y24_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_D = LIOB33_X0Y23_IOB_X0Y23_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_D = LIOB33_X0Y187_IOB_X0Y188_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_D = LIOB33_X0Y187_IOB_X0Y187_I;
  assign LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y208_D = LIOB33_X0Y207_IOB_X0Y208_I;
  assign LIOI3_TBYTESRC_X0Y207_ILOGIC_X0Y207_D = LIOB33_X0Y207_IOB_X0Y207_I;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_A1 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_A2 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_A3 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_A4 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_A5 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_B1 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_B2 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_B3 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_B4 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_B5 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_B6 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_C1 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_C2 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_C3 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_C4 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_C5 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_C6 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_D1 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_D2 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_D3 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_D4 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_D5 = 1'b1;
  assign CLBLL_L_X2Y208_SLICE_X1Y208_D6 = 1'b1;
  assign RIOB33_X105Y95_IOB_X1Y96_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign RIOB33_X105Y95_IOB_X1Y95_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_D4 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_D5 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X72Y145_D6 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A1 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A2 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A4 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A5 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A6 = RIOB33_X105Y155_IOB_X1Y155_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B1 = LIOB33_X0Y17_IOB_X0Y17_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B2 = RIOB33_X105Y157_IOB_X1Y158_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B4 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B5 = LIOB33_X0Y7_IOB_X0Y7_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B6 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C2 = RIOB33_X105Y153_IOB_X1Y154_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C3 = LIOB33_X0Y3_IOB_X0Y4_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C4 = LIOB33_X0Y13_IOB_X0Y13_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C6 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D2 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D3 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D4 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D6 = RIOB33_X105Y155_IOB_X1Y155_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A1 = LIOB33_X0Y3_IOB_X0Y4_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A2 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A3 = LIOB33_X0Y13_IOB_X0Y13_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A4 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A6 = RIOB33_X105Y153_IOB_X1Y154_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B1 = LIOB33_X0Y3_IOB_X0Y4_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B2 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B3 = LIOB33_X0Y13_IOB_X0Y13_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B4 = RIOB33_X105Y153_IOB_X1Y154_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B6 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C2 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C3 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C4 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C6 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D2 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D3 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D4 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D6 = 1'b1;
  assign RIOB33_X105Y97_IOB_X1Y98_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A1 = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A2 = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A3 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A4 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A5 = LIOB33_X0Y241_IOB_X0Y241_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A6 = RIOB33_X105Y151_IOB_X1Y151_I;
  assign RIOB33_X105Y97_IOB_X1Y97_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B3 = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B4 = RIOB33_X105Y151_IOB_X1Y151_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B5 = LIOB33_X0Y241_IOB_X0Y241_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B6 = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C6 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D6 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_R_X59Y159_SLICE_X88Y159_AO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A6 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B6 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C6 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D6 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A1 = LIOB33_X0Y11_IOB_X0Y12_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A2 = LIOB33_X0Y3_IOB_X0Y3_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A3 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A4 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A5 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A6 = RIOB33_X105Y153_IOB_X1Y153_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B1 = CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B2 = CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B3 = CLBLL_L_X2Y102_SLICE_X0Y102_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B4 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B5 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B6 = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_D6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C1 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C2 = LIOB33_X0Y11_IOB_X0Y12_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C3 = LIOB33_X0Y3_IOB_X0Y3_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C4 = RIOB33_X105Y153_IOB_X1Y153_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D6 = 1'b1;
  assign LIOI3_SING_X0Y0_ILOGIC_X0Y0_D = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X44Y158_SLICE_X66Y158_AO5;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A3 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X44Y158_SLICE_X66Y158_BO5;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A6 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_T1 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_D1 = CLBLL_L_X2Y189_SLICE_X0Y189_AO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B1 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B4 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B6 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C2 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C5 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_D1 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C6 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_A1 = LIOB33_X0Y211_IOB_X0Y212_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_A2 = LIOB33_X0Y223_IOB_X0Y224_I;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_T1 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_A4 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_B1 = LIOB33_X0Y211_IOB_X0Y212_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D4 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_T1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D6 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_B2 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_B4 = LIOB33_X0Y235_IOB_X0Y236_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_B5 = LIOB33_X0Y223_IOB_X0Y224_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_B6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_C1 = LIOB33_X0Y215_IOB_X0Y215_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_C2 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_C3 = LIOB33_X0Y239_IOB_X0Y239_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_C4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_C5 = LIOB33_X0Y193_IOB_X0Y193_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_C6 = LIOB33_X0Y227_IOB_X0Y228_I;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_D1 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_D2 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_D3 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_D4 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_D5 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1 = LIOB33_X0Y217_IOB_X0Y217_I;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_A3 = LIOB33_X0Y209_IOB_X0Y210_I;
  assign RIOB33_X105Y101_IOB_X1Y102_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign RIOB33_X105Y101_IOB_X1Y101_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_A5 = LIOB33_X0Y235_IOB_X0Y236_I;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_A1 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_A2 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_A3 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_A6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_A4 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_A5 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_A6 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_B1 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_B2 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_B3 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_B4 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_B5 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_B6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A5 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A6 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_C1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B6 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_C4 = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X44Y158_SLICE_X66Y158_AO5;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X44Y158_SLICE_X66Y158_BO5;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C6 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X0Y210_B3 = LIOB33_X0Y209_IOB_X0Y210_I;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_D1 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_D4 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_D5 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_D6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D6 = 1'b1;
  assign LIOI3_X0Y209_ILOGIC_X0Y210_D = LIOB33_X0Y209_IOB_X0Y210_I;
  assign LIOI3_X0Y209_ILOGIC_X0Y209_D = LIOB33_X0Y209_IOB_X0Y209_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y178_D = LIOB33_X0Y177_IOB_X0Y178_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_D = LIOB33_X0Y177_IOB_X0Y177_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y148_D = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y86_D = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A6 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y85_D = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B6 = 1'b1;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_D = LIOB33_X0Y25_IOB_X0Y26_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_D = LIOB33_X0Y25_IOB_X0Y25_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y214_D = LIOB33_X0Y213_IOB_X0Y214_I;
  assign LIOI3_TBYTETERM_X0Y213_ILOGIC_X0Y213_D = LIOB33_X0Y213_IOB_X0Y213_I;
  assign LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y220_D = LIOB33_X0Y219_IOB_X0Y220_I;
  assign LIOI3_TBYTESRC_X0Y219_ILOGIC_X0Y219_D = LIOB33_X0Y219_IOB_X0Y219_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_D = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_D = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_A6 = CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_A1 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_A2 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_A3 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_A4 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_A5 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_A6 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_B1 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_B2 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_B3 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_B4 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_B5 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_B6 = 1'b1;
  assign RIOB33_X105Y103_IOB_X1Y104_O = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign RIOB33_X105Y103_IOB_X1Y103_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_C1 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_C2 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_C3 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_C4 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_C5 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_C6 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_D1 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_D2 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_D3 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_D4 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_D5 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X67Y152_D6 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_A1 = CLBLM_R_X47Y158_SLICE_X72Y158_BO6;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_A2 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_A3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_A4 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_A5 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_A6 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_B1 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_B2 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_B3 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_B4 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_B5 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_B6 = 1'b1;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X44Y158_SLICE_X66Y158_AO6;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_R_X47Y158_SLICE_X72Y158_AO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_C1 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_C2 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_C3 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_C4 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_C5 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_C6 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_B1 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_D1 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_D2 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_D3 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_D4 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_D5 = 1'b1;
  assign CLBLM_L_X44Y152_SLICE_X66Y152_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_C2 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_C3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_C5 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_C6 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_D2 = 1'b1;
  assign CLBLL_L_X2Y210_SLICE_X1Y210_D3 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1 = 1'b1;
  assign RIOB33_X105Y105_IOB_X1Y106_O = LIOB33_X0Y81_IOB_X0Y81_I;
  assign RIOB33_X105Y105_IOB_X1Y105_O = CLBLL_L_X2Y189_SLICE_X1Y189_AO6;
  assign RIOB33_X105Y165_IOB_X1Y166_O = CLBLM_R_X47Y158_SLICE_X72Y158_AO5;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = LIOB33_X0Y19_IOB_X0Y19_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLL_L_X2Y193_SLICE_X0Y193_AO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = CLBLM_R_X47Y158_SLICE_X72Y158_AO5;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_D1 = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_D1 = CLBLM_L_X44Y158_SLICE_X66Y158_BO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = LIOB33_X0Y19_IOB_X0Y19_I;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = CLBLM_R_X59Y133_SLICE_X88Y133_AO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_D1 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_T1 = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1 = CLBLL_L_X2Y192_SLICE_X0Y192_AO6;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A1 = LIOB33_X0Y1_IOB_X0Y2_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A3 = LIOB33_X0Y243_IOB_X0Y243_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A5 = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A6 = RIOB33_X105Y151_IOB_X1Y152_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C6 = 1'b1;
  assign LIOI3_X0Y241_ILOGIC_X0Y242_D = LIOB33_X0Y241_IOB_X0Y242_I;
  assign LIOI3_X0Y241_ILOGIC_X0Y241_D = LIOB33_X0Y241_IOB_X0Y241_I;
  assign LIOI3_X0Y211_ILOGIC_X0Y212_D = LIOB33_X0Y211_IOB_X0Y212_I;
  assign LIOI3_X0Y211_ILOGIC_X0Y211_D = LIOB33_X0Y211_IOB_X0Y211_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D6 = 1'b1;
  assign LIOI3_X0Y179_ILOGIC_X0Y180_D = LIOB33_X0Y179_IOB_X0Y180_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y179_D = LIOB33_X0Y179_IOB_X0Y179_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_D = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_D = LIOB33_X0Y151_IOB_X0Y151_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_D = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y90_D = LIOB33_X0Y89_IOB_X0Y90_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y89_D = LIOB33_X0Y89_IOB_X0Y89_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A3 = 1'b1;
  assign RIOB33_X105Y107_IOB_X1Y108_O = LIOB33_X0Y201_IOB_X0Y202_I;
  assign RIOB33_X105Y107_IOB_X1Y107_O = LIOB33_X0Y201_IOB_X0Y201_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A6 = 1'b1;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_D = LIOB33_X0Y27_IOB_X0Y28_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B3 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y238_D = LIOB33_X0Y237_IOB_X0Y238_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B4 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y237_ILOGIC_X0Y237_D = LIOB33_X0Y237_IOB_X0Y237_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y232_D = LIOB33_X0Y231_IOB_X0Y232_I;
  assign LIOI3_TBYTESRC_X0Y231_ILOGIC_X0Y231_D = LIOB33_X0Y231_IOB_X0Y231_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_D = LIOB33_X0Y93_IOB_X0Y94_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_D = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D6 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y168_O = LIOB33_X0Y21_IOB_X0Y21_I;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_X0Y19_IOB_X0Y20_I;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_D = RIOB33_X105Y157_IOB_X1Y158_I;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_D = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_C6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A1 = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A2 = LIOB33_X0Y15_IOB_X0Y16_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A3 = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A4 = CLBLL_L_X2Y134_SLICE_X0Y134_BO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A5 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A6 = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B1 = LIOB33_X0Y17_IOB_X0Y18_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B2 = CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B3 = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B4 = LIOB33_X0Y7_IOB_X0Y8_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B5 = RIOB33_X105Y159_IOB_X1Y159_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B6 = LIOB33_X0Y179_IOB_X0Y180_I;
  assign LIOI3_SING_X0Y99_ILOGIC_X0Y99_D = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C1 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C2 = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C4 = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C5 = LIOB33_X0Y15_IOB_X0Y16_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D6 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_A1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_A2 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_A3 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_A4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_A6 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_B1 = CLBLL_L_X2Y189_SLICE_X0Y189_DO6;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_B2 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_B3 = CLBLL_L_X2Y192_SLICE_X0Y192_AO6;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_B4 = CLBLL_L_X2Y194_SLICE_X0Y194_BO6;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_B6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_C1 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_C2 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_C3 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_C4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A1 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X101Y130_D6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A6 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_C5 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_C6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B6 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_D1 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_D2 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X0Y187_D3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D6 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_A1 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_A2 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_A3 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_A4 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_A5 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_A6 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_B1 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_B2 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_B3 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_B4 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_B5 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_B6 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_C1 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_C2 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_C3 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_C4 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_C5 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_C6 = 1'b1;
  assign CLBLM_R_X67Y130_SLICE_X100Y130_A6 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_D1 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_D2 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_D3 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_D4 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_D5 = 1'b1;
  assign CLBLL_L_X2Y187_SLICE_X1Y187_D6 = 1'b1;
  assign RIOB33_X105Y109_IOB_X1Y110_O = LIOB33_X0Y203_IOB_X0Y204_I;
  assign RIOB33_X105Y109_IOB_X1Y109_O = LIOB33_X0Y203_IOB_X0Y203_I;
  assign RIOB33_X105Y169_IOB_X1Y170_O = LIOB33_X0Y23_IOB_X0Y23_I;
  assign RIOB33_X105Y169_IOB_X1Y169_O = LIOB33_X0Y21_IOB_X0Y22_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOB33_X105Y51_IOB_X1Y52_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign RIOB33_X105Y51_IOB_X1Y51_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = LIOB33_X0Y21_IOB_X0Y21_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_D1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_R_X47Y145_SLICE_X73Y145_A4 = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_D1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_T1 = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_D1 = LIOB33_X0Y97_IOB_X0Y97_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_X0Y19_IOB_X0Y20_I;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOB33_X105Y111_IOB_X1Y112_O = CLBLL_L_X2Y192_SLICE_X0Y192_BO6;
  assign RIOB33_X105Y111_IOB_X1Y111_O = LIOB33_X0Y205_IOB_X0Y205_I;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_D1 = CLBLL_L_X2Y189_SLICE_X1Y189_AO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_D1 = CLBLM_L_X44Y152_SLICE_X66Y152_AO6;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1 = CLBLL_L_X2Y193_SLICE_X0Y193_BO6;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = LIOB33_X0Y23_IOB_X0Y23_I;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1 = CLBLL_L_X2Y192_SLICE_X0Y192_BO6;
  assign RIOB33_X105Y171_IOB_X1Y172_O = LIOB33_X0Y25_IOB_X0Y25_I;
  assign RIOB33_X105Y171_IOB_X1Y171_O = LIOB33_X0Y23_IOB_X0Y24_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = LIOB33_X0Y21_IOB_X0Y22_I;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign LIOI3_X0Y215_ILOGIC_X0Y216_D = LIOB33_X0Y215_IOB_X0Y216_I;
  assign LIOI3_X0Y215_ILOGIC_X0Y215_D = LIOB33_X0Y215_IOB_X0Y215_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y184_D = LIOB33_X0Y183_IOB_X0Y184_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y183_D = LIOB33_X0Y183_IOB_X0Y183_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_D = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_D = LIOB33_X0Y153_IOB_X0Y153_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y92_D = LIOB33_X0Y91_IOB_X0Y92_I;
  assign LIOI3_X0Y239_ILOGIC_X0Y240_D = LIOB33_X0Y239_IOB_X0Y240_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y91_D = LIOB33_X0Y91_IOB_X0Y91_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y239_ILOGIC_X0Y239_D = LIOB33_X0Y239_IOB_X0Y239_I;
  assign LIOI3_X0Y1_ILOGIC_X0Y2_D = LIOB33_X0Y1_IOB_X0Y2_I;
  assign LIOI3_X0Y1_ILOGIC_X0Y1_D = LIOB33_X0Y1_IOB_X0Y1_I;
  assign RIOB33_SING_X105Y50_IOB_X1Y50_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_TBYTESRC_X0Y243_ILOGIC_X0Y243_D = LIOB33_X0Y243_IOB_X0Y243_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_A1 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_A2 = LIOB33_X0Y229_IOB_X0Y229_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_A3 = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_A4 = LIOB33_X0Y193_IOB_X0Y194_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_A5 = LIOB33_X0Y215_IOB_X0Y216_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_A6 = CLBLL_L_X2Y187_SLICE_X0Y187_AO5;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_B1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_B2 = LIOB33_X0Y229_IOB_X0Y229_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_B3 = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_B4 = LIOB33_X0Y193_IOB_X0Y194_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_B5 = LIOB33_X0Y215_IOB_X0Y216_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_B6 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_C1 = LIOB33_X0Y233_IOB_X0Y234_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_C2 = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_C3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_C4 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_C5 = LIOB33_X0Y221_IOB_X0Y222_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_C6 = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_D1 = LIOB33_X0Y233_IOB_X0Y234_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_D2 = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_D3 = LIOB33_X0Y221_IOB_X0Y222_I;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_D4 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_D5 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X0Y189_D6 = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign RIOB33_X105Y53_IOB_X1Y53_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOB33_X105Y53_IOB_X1Y54_O = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_A1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_A2 = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_A3 = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_A4 = LIOB33_X0Y221_IOB_X0Y222_I;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_A5 = LIOB33_X0Y233_IOB_X0Y234_I;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_A6 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_SING_X0Y149_ILOGIC_X0Y149_D = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_B1 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_B2 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_B3 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_B4 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_B5 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_B6 = 1'b1;
  assign RIOB33_X105Y113_IOB_X1Y113_O = CLBLL_L_X2Y192_SLICE_X0Y192_BO6;
  assign RIOB33_X105Y113_IOB_X1Y114_O = CLBLL_L_X2Y193_SLICE_X0Y193_BO6;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_C1 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_C2 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_C3 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_C4 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_C5 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_C6 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_D1 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_D2 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_D3 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_D4 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_D5 = 1'b1;
  assign CLBLL_L_X2Y189_SLICE_X1Y189_D6 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = LIOB33_X0Y27_IOB_X0Y28_I;
  assign RIOB33_X105Y173_IOB_X1Y173_O = LIOB33_X0Y27_IOB_X0Y27_I;
  assign RIOB33_SING_X105Y99_IOB_X1Y99_O = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_A1 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_A2 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_A1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_A2 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_A3 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_A6 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_A4 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_A5 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_A6 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_A3 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_B2 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_B3 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_B4 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_B5 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_B6 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_B1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_B2 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_C1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_C1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_C2 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_C3 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_C2 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_C3 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_C4 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_C5 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_C6 = 1'b1;
  assign RIOB33_SING_X105Y100_IOB_X1Y100_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_C4 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_C5 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_C6 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_D1 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_D2 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_D3 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_D4 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_D5 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X89Y159_D6 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_D1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_D2 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X89Y133_D3 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_A2 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_A3 = LIOB33_X0Y239_IOB_X0Y240_I;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_A4 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_A5 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_A6 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_A1 = CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_A2 = CLBLM_R_X47Y158_SLICE_X72Y158_BO6;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_A3 = CLBLL_L_X2Y165_SLICE_X0Y165_BO6;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_A4 = CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_B1 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_B2 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_B3 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_B4 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_B5 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_B6 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_B1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_B2 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_B3 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_B4 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_B5 = 1'b1;
  assign RIOB33_X105Y55_IOB_X1Y56_O = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign RIOB33_X105Y55_IOB_X1Y55_O = CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_B6 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_C1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_C2 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_C3 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_C4 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_C5 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_C6 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_C4 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_C5 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_D1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_D1 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_D2 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_D3 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_D4 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_D5 = 1'b1;
  assign CLBLM_R_X59Y133_SLICE_X88Y133_D6 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_D2 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_D3 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_D4 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_D5 = 1'b1;
  assign CLBLM_R_X59Y159_SLICE_X88Y159_D6 = 1'b1;
  assign RIOB33_X105Y115_IOB_X1Y116_O = CLBLL_L_X2Y192_SLICE_X0Y192_CO6;
  assign RIOB33_X105Y115_IOB_X1Y115_O = CLBLL_L_X2Y193_SLICE_X0Y193_BO6;
endmodule
