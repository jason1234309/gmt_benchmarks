module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y127_IOB_X0Y128_IPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD
  );
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BMUX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CLK;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CLK;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CLK;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CLK;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CLK;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CLK;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5Q;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AQ;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CLK;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BQ;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CLK;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_DO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_DO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CLK;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A5Q;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CLK;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CLK;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CLK;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CLK;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CLK;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CLK;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CLK;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CLK;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5Q;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5Q;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AQ;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CLK;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CLK;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CLK;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CLK;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CQ;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DQ;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CLK;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AQ;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BQ;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CLK;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CQ;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CLK;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AQ;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BQ;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CLK;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BQ;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CLK;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CQ;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CLK;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CLK;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CLK;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CMUX;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AQ;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CLK;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CQ;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DQ;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CLK;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CLK;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CLK;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CLK;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CLK;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CLK;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CLK;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X0Y105_AO5),
.Q(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff0fff0fff0000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc0000aaf0aa33)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_ALUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X1Y105_AO6),
.Q(CLBLL_L_X2Y105_SLICE_X1Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X1Y105_BO6),
.Q(CLBLL_L_X2Y105_SLICE_X1Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000a0f0a000a)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_DLUT (
.I0(CLBLL_L_X2Y105_SLICE_X1Y105_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_CQ),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000010)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_CLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_CQ),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefafafaaeaaaaaa)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_BLUT (
.I0(CLBLL_L_X2Y105_SLICE_X1Y105_DO6),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_CQ),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_DQ),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfccc3000ccff0000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X2Y105_SLICE_X1Y105_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.Q(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.Q(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.Q(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_DO6),
.Q(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hececcecea0a00a0a)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff228822882288)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_CLUT (
.I0(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_DO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa787f7f7f7f)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_DO6),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbfbfbff0f0009c)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_ALUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I3(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000202)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I2(CLBLL_L_X2Y105_SLICE_X1Y105_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000f000e000e000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_ALUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_BO5),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.Q(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000e0e0e020)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_DLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f1fdffffffff)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_CLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc0c0c0ffc060c0)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I2(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.I3(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fbc8f0f0fbfb)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f000f2f2f220)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_DLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.I3(CLBLL_L_X2Y107_SLICE_X1Y107_CO6),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0500cccc05ff)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_CLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafabffbb0000ff33)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0dddf22222222222)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_ALUT (
.I0(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I3(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c14f0f0f050)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_DLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_CO6),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.I4(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.I5(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1450145014500000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_CLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_CO6),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.I4(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4444444444444)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222322255550555)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_ALUT (
.I0(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.Q(CLBLL_L_X2Y108_SLICE_X1Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffeeffceffee)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X0Y108_DO6),
.I1(CLBLL_L_X2Y108_SLICE_X0Y108_CO6),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_DO6),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_CO6),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200323066cc363c)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_CLUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h080a88aaaeafeeff)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_BQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0eac0c0c0eac0c0)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_ALUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I4(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaaffff)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y109_SLICE_X1Y109_AO6),
.Q(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff300030ff030030)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_BQ),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y110_SLICE_X1Y110_BO6),
.Q(CLBLL_L_X2Y110_SLICE_X1Y110_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y110_SLICE_X1Y110_AO6),
.Q(CLBLL_L_X2Y110_SLICE_X1Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aacc0f0f3333)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(CLBLL_L_X2Y110_SLICE_X1Y110_AQ),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_A5Q),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00ff33cc00)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y103_SLICE_X4Y103_AO6),
.Q(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.Q(CLBLL_L_X4Y103_SLICE_X4Y103_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_DO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_CO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf06cf000f000f000)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_BLUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_BQ),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_BO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeccdecc5a005a00)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_ALUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_AQ),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_DO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_CO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_BO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.Q(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000400000000000)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_DLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff80ff)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_CLUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_BQ),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff54ff54ff54)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_BLUT (
.I0(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9d88c888cccc0000)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_BQ),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a000aaaaaaaa)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_ALUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I3(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X4Y105_CO5),
.Q(CLBLL_L_X4Y105_SLICE_X4Y105_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.Q(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0af33333333)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_DLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_BQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_A5Q),
.I4(1'b1),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00003f3faaaa0033)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_CLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_A5Q),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haf00ff00ccdccccc)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_BLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ccccf0e1)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_ALUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I2(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.Q(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddffddffdd55ddff)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_DLUT (
.I0(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I2(1'b1),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I4(CLBLM_R_X5Y106_SLICE_X7Y106_BQ),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080000000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_CLUT (
.I0(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafcfffffafffffff)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I4(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_BQ),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a5a5ff000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_ALUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_DO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I3(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.Q(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.Q(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff1000ffff)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000007fff)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_BQ),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_CQ),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_DO6),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa00fa00ae04ae04)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaabbaab10011001)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_BQ),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.Q(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004550455)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddfffdfffdfffd)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_BQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I3(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ddf5f5ddddf5f5)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_BLUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I4(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000003c003c)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_A5Q),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002000200)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X0Y108_BO6),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010100000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_DO6),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f088f022f022)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff410041ff410041)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.Q(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffffaaaaffff)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcfcfcfcf4)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffef00ef00ef00)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca0cca0cc0acc0a)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.Q(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf555f555ff55ff55)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333337300000050)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.I4(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_BQ),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88d888d888c988c9)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.Q(CLBLL_L_X4Y108_SLICE_X5Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff12ff1200120012)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_A5Q),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc33aa99aaaa)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_C5Q),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000a0a55aa55aa)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_B5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_CQ),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3cff003c3c0000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_DQ),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y103_SLICE_X3Y103_AO6),
.Q(CLBLM_R_X3Y103_SLICE_X3Y103_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff78ff00f0f00000)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_ALUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.I5(CLBLL_L_X4Y103_SLICE_X4Y103_BQ),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.Q(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.Q(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.Q(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffef0f0f0f4f0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I2(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffa5a0e4a0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeefeeddcccdcc)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_CQ),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X3Y104_AO6),
.Q(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.Q(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff5555ffff)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_DLUT (
.I0(CLBLL_L_X4Y103_SLICE_X4Y103_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00003b0800003b08)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_CQ),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffec20cc00)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_BLUT (
.I0(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLL_L_X2Y105_SLICE_X1Y105_BQ),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_CQ),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heccc2000cecc2000)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_ALUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_AQ),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.Q(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.Q(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X2Y105_CO6),
.Q(CLBLM_R_X3Y105_SLICE_X2Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X2Y105_DO6),
.Q(CLBLM_R_X3Y105_SLICE_X2Y105_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafafcf0f0f0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_DLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_CQ),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ddf000f0dd)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_CQ),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf098f01000550055)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_CQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaa00aa00)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0022002233330000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_DLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_CQ),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_DQ),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbeeeebbbbeedd)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_CLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y105_SLICE_X1Y105_BQ),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_DQ),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7d7dbebe)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_BLUT (
.I0(CLBLL_L_X2Y105_SLICE_X1Y105_BQ),
.I1(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y103_SLICE_X4Y103_BQ),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000000080000000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_ALUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_BO5),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_BQ),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_CO6),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_AQ),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_DO6),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.Q(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.Q(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a000000000000)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0707030308080c0c)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_CLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefaaafcccf000)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefceeccfaf0aa00)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.Q(CLBLM_R_X3Y106_SLICE_X3Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.Q(CLBLM_R_X3Y106_SLICE_X3Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.Q(CLBLM_R_X3Y106_SLICE_X3Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf888f888ff888888)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_A5Q),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa0aa0caaa0aa0c)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_CLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_CQ),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f020208888)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_BQ),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'habfa0150aaaa0000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_BQ),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_AQ),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.Q(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLL_L_X2Y107_SLICE_X1Y107_BO6),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfffffffbbff)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_CLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.I1(CLBLL_L_X2Y107_SLICE_X1Y107_BO6),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I5(CLBLL_L_X2Y108_SLICE_X0Y108_BO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0f0e0000000000)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc1100ccfc0030)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_ALUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_CQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_AQ),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.Q(CLBLM_R_X3Y107_SLICE_X3Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.Q(CLBLM_R_X3Y107_SLICE_X3Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0faf0f0f0fef0)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaafffffffbff)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_CLUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5a0a0e4a0e4)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_BQ),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00a0ccccf0f0)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_ALUT (
.I0(CLBLM_R_X3Y107_SLICE_X3Y107_DO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h333300200000ff5f)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.Q(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.Q(CLBLM_R_X3Y108_SLICE_X3Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.Q(CLBLM_R_X3Y108_SLICE_X3Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffbbffbbffbbff)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_CQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd200c3ffe100f0)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_CLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_AO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_CQ),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff90ff9090909090)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_BLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_BQ),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.I3(CLBLM_R_X3Y108_SLICE_X3Y108_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hecdcecdca050a050)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_ALUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.I1(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.I3(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_BO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_DO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffecececffa0a0a0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_CQ),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_DQ),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff888f888f888)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_CQ),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefaaafcccf000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefceeccfaf0aa00)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.Q(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00ff00)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_BO6),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fcf3fcf3fcf3ed)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_BQ),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_CQ),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_DQ),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ff6ffffffff6ff6)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_DQ),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_CQ),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_AQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccbf00cccc4000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_BQ),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.Q(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.Q(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200ffffddffddff)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_CLUT (
.I0(CLBLM_R_X5Y104_SLICE_X7Y104_DQ),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haac0aac0aa30aa30)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_BLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22cc00dc10dc10)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y104_SLICE_X7Y104_AO6),
.Q(CLBLM_R_X5Y104_SLICE_X7Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y104_SLICE_X7Y104_BO6),
.Q(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y104_SLICE_X7Y104_CO6),
.Q(CLBLM_R_X5Y104_SLICE_X7Y104_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y104_SLICE_X7Y104_DO6),
.Q(CLBLM_R_X5Y104_SLICE_X7Y104_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd88c8888d8d88888)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X5Y104_SLICE_X7Y104_CQ),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_DQ),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc0100000c0c0)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_CLUT (
.I0(CLBLM_R_X5Y104_SLICE_X7Y104_DQ),
.I1(CLBLM_R_X5Y104_SLICE_X7Y104_CQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f020f088f020)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00a0a00202)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_AQ),
.I3(CLBLM_R_X5Y104_SLICE_X7Y104_DQ),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.Q(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.Q(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X6Y105_CO6),
.Q(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccecccccccccc8)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_DLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_AQ),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_CQ),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000009888)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f044440014)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff40ff4100400041)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_CQ),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.Q(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.Q(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.Q(CLBLM_R_X5Y105_SLICE_X7Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_DLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_CQ),
.I2(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.I4(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff005808f000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_CLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_CO5),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_CQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc58cc88cc08cc88)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_CO5),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc10dc10dc01dc01)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8c008c00bf33bf33)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_DLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_BQ),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff02ff02ff)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002330000)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I5(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafaaaeafaf)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_ALUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.I4(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I5(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.Q(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.Q(CLBLM_R_X5Y106_SLICE_X7Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0c030c03)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_BLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000062aa4000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_CO5),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.Q(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000008880000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff755ffff)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_DO6),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccccc4ccc)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_BLUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_BQ),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfc0030cccf0003)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.Q(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffff0f0f0f0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_CLUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_BQ),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffddfdddffdd)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_BLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I1(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa31aa33aa02aa00)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_ALUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_BQ),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.Q(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.Q(CLBLM_R_X5Y108_SLICE_X6Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffffffffffffff)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_DLUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_AQ),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_CQ),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888fff7ffff)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_CLUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_BQ),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf09cf0ccf000f000)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_BLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_BQ),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hebaa5000ebaa5000)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.Q(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.Q(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.Q(CLBLM_R_X5Y108_SLICE_X7Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7fffff7f7f)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_DLUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_CQ),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8f2f808080808)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_CQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_AQ),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4b1a0a0e4b1)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BQ),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_CQ),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa05aa00fa50aa00)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_AQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X3Y107_AQ),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X1Y108_AQ),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X1Y108_AQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y128_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D = CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_BMUX = CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A = CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_AMUX = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_BMUX = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_AMUX = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_AMUX = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_BMUX = CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_AMUX = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_BMUX = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_BMUX = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_CMUX = CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_AMUX = CLBLL_L_X2Y110_SLICE_X1Y110_A5Q;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_BMUX = CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A = CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D = CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_AMUX = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_AMUX = CLBLL_L_X4Y105_SLICE_X4Y105_A5Q;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_BMUX = CLBLL_L_X4Y105_SLICE_X4Y105_BO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_CMUX = CLBLL_L_X4Y105_SLICE_X4Y105_CO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_DMUX = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_CMUX = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_BMUX = CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_BMUX = CLBLL_L_X4Y109_SLICE_X4Y109_B5Q;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_CMUX = CLBLL_L_X4Y109_SLICE_X4Y109_C5Q;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C = CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D = CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_AMUX = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_BMUX = CLBLM_R_X3Y105_SLICE_X2Y105_BO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_CMUX = CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_AMUX = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_CMUX = CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C = CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D = CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_CMUX = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_CMUX = CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_DMUX = CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_R_X3Y107_SLICE_X3Y107_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C3 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C4 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A2 = CLBLM_R_X3Y106_SLICE_X3Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A3 = CLBLM_R_X3Y106_SLICE_X3Y106_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A4 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A5 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B2 = CLBLM_R_X3Y106_SLICE_X3Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B3 = CLBLM_R_X3Y106_SLICE_X3Y106_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B5 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C1 = CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C2 = CLBLM_R_X3Y106_SLICE_X3Y106_CQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D2 = CLBLL_L_X4Y105_SLICE_X4Y105_A5Q;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D3 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D4 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D5 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D6 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A3 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A4 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A5 = CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B2 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B3 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B5 = CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C1 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C5 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D1 = CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D5 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D6 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_R_X3Y107_SLICE_X3Y107_AQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A2 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A3 = CLBLM_R_X5Y104_SLICE_X7Y104_AQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A4 = CLBLM_R_X5Y104_SLICE_X7Y104_DQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A5 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B2 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B3 = CLBLM_R_X5Y104_SLICE_X7Y104_AQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B5 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B6 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A1 = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A2 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A4 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A6 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C1 = CLBLM_R_X5Y104_SLICE_X7Y104_DQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C2 = CLBLM_R_X5Y104_SLICE_X7Y104_CQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B2 = CLBLM_R_X3Y107_SLICE_X3Y107_BQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B3 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B5 = CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C1 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C2 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C3 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C4 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C5 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C6 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D2 = CLBLM_R_X5Y104_SLICE_X7Y104_CQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D3 = CLBLM_R_X5Y104_SLICE_X7Y104_DQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A4 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A3 = CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D1 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D2 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D3 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D4 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A6 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B1 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B2 = CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A1 = CLBLM_R_X3Y106_SLICE_X3Y106_CQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A3 = CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A5 = CLBLM_R_X3Y107_SLICE_X3Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B6 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C1 = CLBLM_R_X5Y104_SLICE_X7Y104_DQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C2 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B2 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B3 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B4 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B5 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B6 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D2 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C1 = CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C2 = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C3 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C4 = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C5 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C6 = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D4 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C6 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D2 = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D3 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D4 = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D5 = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D6 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A3 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A4 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A6 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B2 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B3 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B5 = CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B6 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B4 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B5 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A1 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A2 = CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A3 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A4 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C1 = CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C2 = CLBLM_R_X5Y105_SLICE_X7Y105_CQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B1 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B2 = CLBLM_R_X3Y108_SLICE_X3Y108_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B3 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B4 = CLBLM_R_X3Y108_SLICE_X3Y108_CQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D1 = CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D2 = CLBLM_R_X5Y105_SLICE_X7Y105_CQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C1 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C2 = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C3 = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C5 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C6 = CLBLM_R_X3Y108_SLICE_X3Y108_CQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D3 = CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D4 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A2 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A3 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A5 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D1 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D2 = CLBLM_R_X3Y108_SLICE_X3Y108_CQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D4 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A6 = CLBLM_R_X5Y105_SLICE_X7Y105_CQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B2 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B3 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B4 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A3 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A5 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C1 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C2 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B5 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B6 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D1 = CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D2 = CLBLL_L_X2Y110_SLICE_X1Y110_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D3 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D4 = CLBLM_R_X5Y105_SLICE_X7Y105_CQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D6 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C5 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C6 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A2 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A3 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A4 = CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A5 = CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B1 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B2 = CLBLM_R_X5Y106_SLICE_X7Y106_BQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B4 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = CLBLM_R_X3Y108_SLICE_X3Y108_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = CLBLM_R_X3Y109_SLICE_X2Y109_DQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = CLBLM_R_X3Y108_SLICE_X3Y108_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = CLBLL_L_X4Y109_SLICE_X4Y109_CQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = CLBLM_R_X3Y108_SLICE_X3Y108_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = CLBLM_R_X3Y109_SLICE_X2Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = CLBLM_R_X3Y109_SLICE_X2Y109_DQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = CLBLL_L_X4Y109_SLICE_X4Y109_B5Q;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A1 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A2 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A3 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A4 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A5 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A6 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B1 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B2 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B3 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B6 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C1 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C2 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C6 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D1 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D2 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = CLBLM_R_X3Y109_SLICE_X2Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D3 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D4 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D6 = CLBLM_R_X5Y106_SLICE_X7Y106_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = CLBLM_R_X3Y109_SLICE_X2Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = CLBLM_R_X3Y109_SLICE_X2Y109_DQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A1 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A2 = CLBLL_L_X2Y105_SLICE_X1Y105_AQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A3 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A4 = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B1 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B2 = CLBLL_L_X4Y103_SLICE_X4Y103_BQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B3 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B6 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C1 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C2 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C4 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D1 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D2 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D4 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A1 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A2 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A4 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B1 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B2 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B4 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A1 = CLBLM_R_X5Y108_SLICE_X6Y108_BQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A3 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C1 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C2 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C4 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A5 = CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A6 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B1 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B2 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B3 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B4 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B5 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D1 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D2 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D4 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C1 = CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C2 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C3 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C4 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C5 = CLBLM_R_X5Y108_SLICE_X6Y108_BQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C6 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D4 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A3 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A5 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A6 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B1 = CLBLM_R_X5Y108_SLICE_X6Y108_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B3 = CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B4 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B5 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B6 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C1 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C2 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C3 = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C4 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C5 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C6 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D1 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D2 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D3 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D4 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D5 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D6 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C4 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C6 = CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D4 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D6 = CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A2 = CLBLM_R_X3Y106_SLICE_X3Y106_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A3 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A5 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B1 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B2 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B3 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B4 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B5 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B6 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C1 = CLBLM_R_X3Y106_SLICE_X3Y106_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C2 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C3 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C4 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C5 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C6 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D1 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D2 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D3 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D4 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D6 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A1 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A2 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A3 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A4 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A5 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A6 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B1 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B2 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B3 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B4 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C1 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C2 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C3 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C4 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A3 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A4 = CLBLL_L_X4Y108_SLICE_X5Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A6 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B2 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D1 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D2 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D3 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D4 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C2 = CLBLM_R_X5Y108_SLICE_X7Y108_CQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C4 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C5 = CLBLL_L_X4Y108_SLICE_X5Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C6 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D1 = CLBLM_R_X5Y108_SLICE_X7Y108_CQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D2 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D3 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D4 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D5 = CLBLL_L_X4Y108_SLICE_X5Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C4 = CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A2 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A3 = CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A5 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C5 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B1 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B2 = CLBLM_R_X5Y108_SLICE_X6Y108_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B3 = CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B5 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C1 = CLBLM_R_X5Y108_SLICE_X6Y108_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C2 = CLBLM_R_X5Y108_SLICE_X6Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C3 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C4 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C5 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D1 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D2 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D3 = CLBLL_L_X4Y108_SLICE_X5Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D4 = CLBLM_R_X5Y108_SLICE_X7Y108_CQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D5 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D6 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A1 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A2 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A3 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A4 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_AX = CLBLL_L_X4Y105_SLICE_X4Y105_CO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B1 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B3 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B4 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B5 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C1 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C4 = CLBLL_L_X4Y105_SLICE_X4Y105_A5Q;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D1 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D2 = CLBLM_R_X5Y106_SLICE_X7Y106_BQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D3 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D4 = CLBLL_L_X4Y105_SLICE_X4Y105_A5Q;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D6 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A1 = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A3 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A4 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B1 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B2 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B3 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B4 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B5 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B6 = CLBLM_R_X5Y106_SLICE_X7Y106_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C1 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C2 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C3 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C4 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C5 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C6 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D1 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D2 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D4 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D5 = CLBLM_R_X5Y106_SLICE_X7Y106_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B6 = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A3 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A4 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A6 = CLBLM_R_X5Y106_SLICE_X7Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B2 = CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B4 = CLBLM_R_X3Y107_SLICE_X3Y107_BQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A1 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A2 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A3 = CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C2 = CLBLM_R_X3Y106_SLICE_X3Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C3 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B3 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B5 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C4 = CLBLM_R_X3Y106_SLICE_X3Y106_CQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C5 = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D1 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D2 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D3 = CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D4 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D5 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D6 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A2 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A3 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A5 = CLBLL_L_X4Y105_SLICE_X4Y105_A5Q;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B1 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B3 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B4 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A3 = CLBLL_L_X2Y105_SLICE_X1Y105_AQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A4 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A5 = CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C1 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C2 = CLBLM_R_X5Y106_SLICE_X7Y106_BQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B1 = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B2 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B4 = CLBLM_R_X3Y105_SLICE_X2Y105_CQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B6 = CLBLM_R_X3Y105_SLICE_X2Y105_DQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C3 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C4 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C1 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C2 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C5 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C6 = CLBLM_R_X3Y105_SLICE_X2Y105_CQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D6 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D1 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D2 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D3 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D4 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D1 = CLBLL_L_X2Y105_SLICE_X1Y105_BQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D4 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D6 = CLBLM_R_X3Y105_SLICE_X2Y105_CQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A1 = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A2 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A3 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A4 = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_AX = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B1 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B2 = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B3 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C1 = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C2 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C4 = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C6 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D2 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D3 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D5 = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A1 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A2 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A3 = CLBLM_R_X3Y105_SLICE_X2Y105_BO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A4 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A6 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B2 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B3 = CLBLL_L_X2Y105_SLICE_X1Y105_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B6 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_R_X3Y107_SLICE_X3Y107_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A2 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A3 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A4 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A5 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = CLBLM_R_X5Y108_SLICE_X7Y108_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = CLBLM_R_X3Y107_SLICE_X3Y107_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B1 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B2 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B3 = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B4 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B6 = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C1 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C2 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C3 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C4 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C6 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D2 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D3 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D4 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D6 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = CLBLL_L_X4Y108_SLICE_X5Y108_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = CLBLL_L_X2Y110_SLICE_X1Y110_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A1 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A3 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A4 = CLBLM_R_X3Y108_SLICE_X3Y108_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A5 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B1 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B3 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B5 = CLBLM_R_X3Y108_SLICE_X3Y108_CQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C1 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C4 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C5 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C6 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D2 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D3 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D4 = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D5 = CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D6 = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C4 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C5 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = CLBLM_R_X3Y109_SLICE_X2Y109_DQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D5 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = CLBLL_L_X4Y109_SLICE_X4Y109_B5Q;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = CLBLL_L_X4Y109_SLICE_X4Y109_CQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A1 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A3 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = CLBLL_L_X4Y109_SLICE_X4Y109_C5Q;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_C5Q;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B3 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B5 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C1 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C2 = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C3 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C4 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C5 = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C6 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D2 = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D3 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D4 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D5 = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D6 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A1 = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A3 = CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A4 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A5 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B1 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B3 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B4 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B5 = CLBLM_R_X3Y108_SLICE_X3Y108_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C1 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C2 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C3 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C4 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D2 = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D3 = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D4 = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D5 = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D6 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B5 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A1 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A2 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A3 = CLBLM_R_X3Y103_SLICE_X3Y103_AQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A5 = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A6 = CLBLL_L_X4Y103_SLICE_X4Y103_BQ;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B6 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C6 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C3 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C4 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B6 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C6 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = CLBLM_R_X3Y108_SLICE_X3Y108_BQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A1 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A3 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A5 = CLBLM_R_X3Y103_SLICE_X3Y103_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A6 = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B1 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B4 = CLBLL_L_X2Y105_SLICE_X1Y105_BQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B5 = CLBLM_R_X3Y105_SLICE_X2Y105_CQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B6 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C2 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C3 = CLBLM_R_X3Y105_SLICE_X2Y105_CQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C4 = CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D1 = CLBLL_L_X4Y103_SLICE_X4Y103_BQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D5 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A2 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A3 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A6 = CLBLM_R_X3Y106_SLICE_X3Y106_CQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A4 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B3 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B4 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B6 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C2 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C3 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C4 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C6 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B3 = CLBLM_R_X5Y108_SLICE_X7Y108_CQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B4 = CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B5 = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_BX = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_AX = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = CLBLL_L_X2Y110_SLICE_X1Y110_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = CLBLL_L_X2Y110_SLICE_X1Y110_A5Q;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A1 = CLBLL_L_X4Y105_SLICE_X4Y105_BO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A2 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A3 = CLBLL_L_X4Y103_SLICE_X4Y103_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A4 = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A5 = CLBLM_R_X3Y103_SLICE_X3Y103_AQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A6 = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B1 = CLBLL_L_X2Y105_SLICE_X1Y105_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B2 = CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B3 = CLBLM_R_X3Y103_SLICE_X3Y103_AQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B5 = CLBLL_L_X4Y103_SLICE_X4Y103_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B6 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C1 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C2 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C4 = CLBLL_L_X2Y105_SLICE_X1Y105_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C5 = CLBLM_R_X3Y105_SLICE_X2Y105_DQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C6 = CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D4 = CLBLM_R_X3Y105_SLICE_X2Y105_CQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D5 = CLBLM_R_X3Y105_SLICE_X2Y105_DQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D6 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A2 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_AX = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B2 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B3 = CLBLM_R_X3Y105_SLICE_X2Y105_CQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B5 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C1 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C2 = CLBLM_R_X3Y105_SLICE_X2Y105_CQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C3 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D2 = CLBLM_R_X3Y105_SLICE_X2Y105_CQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D3 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D4 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C1 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
endmodule
