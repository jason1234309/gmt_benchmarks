module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y63_IOB_X0Y64_OPAD,
  output LIOB33_X0Y65_IOB_X0Y65_OPAD,
  output LIOB33_X0Y65_IOB_X0Y66_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_AO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_AO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_BO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_BO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_CO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_CO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_DO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_DO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_AO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_AO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_BO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_BO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_BQ;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_CLK;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_CO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_CO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_DO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_DO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_DQ;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_AMUX;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_AO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_AO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_AQ;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_BO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_CLK;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_CO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_CO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_DO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_DO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_AO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_AO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_AQ;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_BO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_BO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C5Q;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_CLK;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_CMUX;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_CO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_CO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_CQ;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_DO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_DO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AQ;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BQ;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CLK;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_DO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_DO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_AO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_AO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_AQ;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B5Q;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BQ;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_CLK;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_CO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_CO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_DO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_DO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_AO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_AO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_BO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_BO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_BQ;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CLK;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CQ;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_DO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_DO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_DQ;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_AO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_BO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_BO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_CO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_CO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_DO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_DO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_AO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_AO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_BO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_BO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_CO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_CO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_DO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_DO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CMUX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DMUX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C5Q;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CLK;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CLK;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D5Q;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CLK;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CLK;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CLK;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CLK;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CLK;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CLK;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CLK;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CLK;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CLK;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CLK;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CE;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CLK;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C5Q;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CLK;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AMUX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C5Q;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CLK;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CMUX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C5Q;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CLK;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CMUX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DMUX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C5Q;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CLK;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A5Q;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C5Q;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CLK;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C5Q;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CLK;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CLK;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CMUX;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A5Q;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AMUX;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DMUX;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B5Q;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CLK;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C5Q;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CLK;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CLK;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CE;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CLK;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A5Q;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CLK;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B5Q;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BMUX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C5Q;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CLK;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CMUX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CE;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CLK;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CE;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CLK;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_DO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C5Q;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CLK;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CLK;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CE;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CLK;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CLK;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CLK;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CLK;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CLK;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AMUX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_DO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_DO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_DO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_DO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_DO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_AMUX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_AO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_BMUX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_BO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CMUX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_DO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_DO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AMUX;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5Q;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5Q;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A5Q;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CE;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B5Q;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CLK;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CLK;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CE;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CLK;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CLK;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CLK;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CLK;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CE;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CLK;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CLK;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_DO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B5Q;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C5Q;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D5Q;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B5Q;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CLK;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C5Q;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CLK;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A5Q;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AMUX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BMUX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CLK;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AMUX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BMUX;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CLK;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AMUX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AMUX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AMUX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BMUX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CLK;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BMUX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AMUX;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AMUX;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CLK;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AMUX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BMUX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CE;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CLK;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DMUX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CLK;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BMUX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CLK;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CLK;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_AMUX;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_AO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_AO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_BMUX;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_BO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_CMUX;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_CO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_CO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_DO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_DO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_BO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_CO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_CO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_DO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A5Q;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AMUX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BMUX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CLK;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CLK;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A5Q;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CLK;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B5Q;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C5Q;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CLK;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CLK;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A5Q;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AMUX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_BO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_BO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CLK;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_DO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_DO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_DQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C5Q;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CLK;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CMUX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D5Q;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DMUX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AMUX;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AX;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BMUX;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BX;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CE;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CLK;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_DO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_DO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C5Q;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CLK;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CMUX;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_DO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_DO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CLK;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_DMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_DO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_DO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A5Q;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B5Q;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CLK;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D5Q;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CLK;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D5Q;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B5Q;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C5Q;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CLK;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A5Q;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AMUX;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CLK;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AMUX;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B5Q;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BMUX;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C5Q;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CLK;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CMUX;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D5Q;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DMUX;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AMUX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BMUX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CE;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CLK;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CMUX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DMUX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AMUX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B5Q;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BMUX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C5Q;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CLK;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CMUX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_DO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A5Q;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AMUX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_BO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_BO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_BQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CLK;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CMUX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_DO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AMUX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CLK;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CMUX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DMUX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CLK;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CLK;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CLK;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_A;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_A1;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_A2;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_A3;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_A4;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_A5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_A6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_AO5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_AO6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_A_CY;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_A_XOR;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_B;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_B1;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_B2;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_B3;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_B4;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_B5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_B6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_BO5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_BO6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_B_CY;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_B_XOR;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_C;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_C1;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_C2;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_C3;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_C4;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_C5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_C6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_CO5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_CO6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_C_CY;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_C_XOR;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_D;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_D1;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_D2;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_D3;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_D4;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_D5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_D6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_DO5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_DO6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_D_CY;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X2Y165_D_XOR;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_A;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_A1;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_A2;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_A3;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_A4;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_A5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_A6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_AO5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_AO6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_A_CY;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_A_XOR;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_B;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_B1;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_B2;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_B3;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_B4;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_B5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_B6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_BO5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_BO6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_B_CY;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_B_XOR;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_C;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_C1;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_C2;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_C3;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_C4;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_C5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_C6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_CO5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_CO6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_C_CY;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_C_XOR;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_D;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_D1;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_D2;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_D3;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_D4;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_D5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_D6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_DO5;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_DO6;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_D_CY;
  wire [0:0] CLBLM_R_X3Y165_SLICE_X3Y165_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C5Q;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CLK;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CLK;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CLK;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D5Q;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A5Q;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B5Q;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C5Q;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CLK;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B5Q;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C5Q;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CLK;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D5Q;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CLK;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_DO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C5Q;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CLK;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A5Q;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B5Q;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C5Q;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CLK;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A5Q;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AMUX;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CLK;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A5Q;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AMUX;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CLK;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CLK;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CLK;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B5Q;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C5Q;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A5Q;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CLK;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B5Q;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CLK;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CLK;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CE;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CLK;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CLK;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B5Q;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CLK;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C5Q;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CLK;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B5Q;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C5Q;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CLK;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A5Q;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CLK;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A5Q;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CLK;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CLK;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CE;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CLK;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CLK;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B5Q;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CLK;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D5Q;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C5Q;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CLK;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C5Q;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D5Q;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A5Q;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_O;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_TQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_TQ;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_DO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_CO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_BO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y55_IOB_X0Y56_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_AO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_DO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_CO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_BO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_AO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_DO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_CO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_BO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_AO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y135_SLICE_X1Y135_AO6),
.Q(CLBLL_L_X2Y135_SLICE_X1Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y135_SLICE_X1Y135_BO6),
.Q(CLBLL_L_X2Y135_SLICE_X1Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y135_SLICE_X1Y135_CO6),
.Q(CLBLL_L_X2Y135_SLICE_X1Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y135_SLICE_X1Y135_DO6),
.Q(CLBLL_L_X2Y135_SLICE_X1Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaf0005aafa0050)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLL_L_X2Y135_SLICE_X1Y135_DQ),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_DQ),
.I4(CLBLL_L_X2Y135_SLICE_X1Y135_AQ),
.I5(CLBLM_R_X3Y135_SLICE_X2Y135_BO6),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_DO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888888d8d8)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_C5Q),
.I2(CLBLL_L_X2Y135_SLICE_X1Y135_BQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y135_SLICE_X1Y135_AQ),
.I5(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_CO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888d88dd8888)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y138_SLICE_X1Y138_BQ),
.I2(CLBLL_L_X2Y135_SLICE_X1Y135_AQ),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I5(CLBLL_L_X2Y135_SLICE_X1Y135_BQ),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_BO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000caaaa00f0)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I2(CLBLL_L_X2Y135_SLICE_X1Y135_AQ),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X2Y135_SLICE_X1Y135_BQ),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_AO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y137_SLICE_X0Y137_AO6),
.Q(CLBLL_L_X2Y137_SLICE_X0Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X0Y137_DO5),
.O6(CLBLL_L_X2Y137_SLICE_X0Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X0Y137_CO5),
.O6(CLBLL_L_X2Y137_SLICE_X0Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X0Y137_BO5),
.O6(CLBLL_L_X2Y137_SLICE_X0Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc5accf00000ffff)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_ALUT (
.I0(CLBLM_R_X3Y138_SLICE_X2Y138_DQ),
.I1(CLBLM_R_X3Y137_SLICE_X2Y137_D5Q),
.I2(CLBLL_L_X2Y137_SLICE_X0Y137_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(LIOB33_X0Y59_IOB_X0Y60_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X0Y137_AO5),
.O6(CLBLL_L_X2Y137_SLICE_X0Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y137_SLICE_X1Y137_CO5),
.Q(CLBLL_L_X2Y137_SLICE_X1Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y137_SLICE_X1Y137_AO6),
.Q(CLBLL_L_X2Y137_SLICE_X1Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y137_SLICE_X1Y137_BO6),
.Q(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y137_SLICE_X1Y137_CO6),
.Q(CLBLL_L_X2Y137_SLICE_X1Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X1Y137_DO5),
.O6(CLBLL_L_X2Y137_SLICE_X1Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaccccf0f0)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_CLUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I1(CLBLL_L_X2Y137_SLICE_X1Y137_CQ),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X1Y137_CO5),
.O6(CLBLL_L_X2Y137_SLICE_X1Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff88ffaa008800aa)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_BLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I1(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.O5(CLBLL_L_X2Y137_SLICE_X1Y137_BO5),
.O6(CLBLL_L_X2Y137_SLICE_X1Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafff03330)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_ALUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_DQ),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I2(CLBLL_L_X2Y137_SLICE_X1Y137_AQ),
.I3(CLBLL_L_X2Y137_SLICE_X1Y137_CQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X2Y137_SLICE_X1Y137_AO5),
.O6(CLBLL_L_X2Y137_SLICE_X1Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_DO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_CO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_BO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_AO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y138_SLICE_X1Y138_AO6),
.Q(CLBLL_L_X2Y138_SLICE_X1Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y138_SLICE_X1Y138_BO6),
.Q(CLBLL_L_X2Y138_SLICE_X1Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_DO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_CO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeeeaaaa14440000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y138_SLICE_X1Y138_BQ),
.I2(CLBLL_L_X2Y138_SLICE_X1Y138_AQ),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_CO6),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I5(CLBLM_R_X3Y138_SLICE_X3Y138_B5Q),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_BO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3c00aaaa3c00)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_ALUT (
.I0(CLBLL_L_X2Y139_SLICE_X0Y139_B5Q),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_CO6),
.I2(CLBLL_L_X2Y138_SLICE_X1Y138_AQ),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_AO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y139_SLICE_X0Y139_BO5),
.Q(CLBLL_L_X2Y139_SLICE_X0Y139_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y139_SLICE_X0Y139_AO6),
.Q(CLBLL_L_X2Y139_SLICE_X0Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y139_SLICE_X0Y139_BO6),
.Q(CLBLL_L_X2Y139_SLICE_X0Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_DO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_CO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaccaacc)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_BLUT (
.I0(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_C5Q),
.I2(CLBLL_L_X2Y139_SLICE_X0Y139_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_BO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2f3f3e2e2f3f3)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_AO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y139_SLICE_X1Y139_AO6),
.Q(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y139_SLICE_X1Y139_BO6),
.Q(CLBLL_L_X2Y139_SLICE_X1Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y139_SLICE_X1Y139_CO6),
.Q(CLBLL_L_X2Y139_SLICE_X1Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y139_SLICE_X1Y139_DO6),
.Q(CLBLL_L_X2Y139_SLICE_X1Y139_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d888d88d888d888)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.I2(CLBLL_L_X2Y139_SLICE_X1Y139_DQ),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y139_SLICE_X2Y139_CO6),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_DO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf00c00f6f00600)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_CLUT (
.I0(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I1(CLBLL_L_X2Y139_SLICE_X1Y139_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.I5(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_CO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f08800f0f0aa00)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_BLUT (
.I0(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.I1(CLBLL_L_X2Y139_SLICE_X1Y139_BQ),
.I2(CLBLL_L_X2Y137_SLICE_X1Y137_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y139_SLICE_X2Y139_BO6),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_BO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0caaccaaccaacc)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_ALUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I1(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.I2(CLBLM_R_X3Y138_SLICE_X2Y138_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y137_SLICE_X0Y137_AQ),
.I5(LIOB33_X0Y59_IOB_X0Y60_I),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_AO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_AO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_DLUT (
.I0(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I5(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000080000000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_CLUT (
.I0(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hba10ba10ea40ea40)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I2(LIOB33_X0Y53_IOB_X0Y54_I),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_CO6),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf15bf15fb51fb51)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y129_SLICE_X3Y129_BO5),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_AO6),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_BO6),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_CO6),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f00000f0f0000)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_DO6),
.I3(1'b1),
.I4(LIOB33_X0Y53_IOB_X0Y54_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fcf0f0030c0000)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff002828ff002828)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_BLUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_CO5),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7df500007df5)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_ALUT (
.I0(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_AO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_DO5),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_CO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc000000a3afaca0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_DLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3aca3accfcfc0c0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_CLUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaa400000ff00ff)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55bb11fa50ba10)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I3(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I5(CLBLM_R_X3Y133_SLICE_X2Y133_CQ),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_CO5),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_DO5),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_AO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_BO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_CO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_DO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ffcc00cc)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y133_SLICE_X5Y133_C5Q),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccff00)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fa50ee44)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_C5Q),
.I3(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I4(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaafefe54005454)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I5(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_BO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_CO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a000a000a000)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0bbbbeeee)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I2(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q),
.I3(1'b1),
.I4(CLBLL_L_X4Y132_SLICE_X4Y132_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb88bb88bb)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_BLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_A5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y134_SLICE_X5Y134_CO6),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe3232ccfe0032)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_ALUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_AO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_BO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_CLUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_DO6),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I5(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5ccffccfaccf0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_C5Q),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaac0aaffaacc)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_DO6),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_CO6),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_CO5),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_DO5),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_CO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_DO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0aaf0aaf0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_DLUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_C5Q),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0f0aaf0aa)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_CLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa0fccaaccaa)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_BLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_CQ),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbb00bbffb000b0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_C5Q),
.I5(CLBLM_R_X3Y133_SLICE_X2Y133_C5Q),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_CO5),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_AO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_CO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffefffe)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_DLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfa0afa0a)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_CLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_D5Q),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff003030fcfc)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb888b8bbb888b8)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_ALUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_BO5),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_AO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_BO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7080000ff000000)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_DLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_DO6),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I4(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff3fff3fff)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1d1d1d1fc30fc30)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_BLUT (
.I0(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ff00fafa)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_ALUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_DO6),
.I1(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff5fffffffff)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_BO5),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7ffffffffff)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_BO5),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffc7f7f7f7f)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_BLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffccffcc)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y133_SLICE_X5Y133_DO6),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.I3(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_AO5),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_BO5),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_DO5),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_AO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_BO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_CO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_DO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d8d8d8dee44ee44)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_DO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffef5545ffff5555)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I5(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_CO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0bbbb8888)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_BLUT (
.I0(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_BO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ffcccc00ff)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_ALUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_DQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_C5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_AO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_AO5),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_AO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ff66ffff66ff66)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_DLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_D5Q),
.I1(CLBLL_L_X2Y138_SLICE_X1Y138_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_B5Q),
.I4(1'b1),
.I5(CLBLL_L_X2Y138_SLICE_X1Y138_BQ),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_DO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d7dbebe7d7dbebe)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_CLUT (
.I0(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_BQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_CO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7bffdeff)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_BLUT (
.I0(CLBLM_R_X3Y137_SLICE_X2Y137_DQ),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I2(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.I4(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I5(CLBLL_L_X4Y135_SLICE_X5Y135_CO6),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_BO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaaaffaa00)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_ALUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_AO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_AO5),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_BO5),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_CO5),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_DO5),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_AO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_BO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_CO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_DO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccff3c003c)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_DLUT (
.I0(CLBLL_L_X2Y138_SLICE_X1Y138_AQ),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_DO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88f3f3c0c0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_CLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I3(CLBLL_L_X4Y131_SLICE_X5Y131_D5Q),
.I4(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_CO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222f3c0f3c0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y122_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_B5Q),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_BO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f000ff0ccf0cc)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_AO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_CO5),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_AO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_DO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffaaf0f05500)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_A5Q),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_DO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbebe1414ff55aa00)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_DO6),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_CO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cfcff000ff0f)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22fc30ee22ee22)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I3(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_AO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_CO5),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_DO5),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_CO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_DO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f000ccf0ccf0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_DLUT (
.I0(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_DO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc33008bb88bb8)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_CLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y137_SLICE_X2Y137_D5Q),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_CO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff44f0f0bb00)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_BLUT (
.I0(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I1(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_DQ),
.I3(CLBLM_R_X3Y138_SLICE_X2Y138_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_BO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aae2aae2)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_ALUT (
.I0(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_CO5),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_DO5),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_AO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_BO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_CO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_DO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222f3c0f3c0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y137_SLICE_X5Y137_DQ),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_DO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5a0f5a0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_D5Q),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_C5Q),
.I3(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_CO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000003f)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_BLUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_B5Q),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.I2(CLBLL_L_X4Y137_SLICE_X5Y137_AQ),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_DQ),
.I4(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_BO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffffffcc)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_ALUT (
.I0(CLBLM_R_X3Y133_SLICE_X2Y133_B5Q),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_DQ),
.I4(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_AO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_CQ),
.Q(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfc)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_CQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y138_SLICE_X8Y138_A5Q),
.I5(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000000)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_CLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_C5Q),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I3(1'b1),
.I4(CLBLL_L_X4Y138_SLICE_X4Y138_DO6),
.I5(CLBLL_L_X4Y138_SLICE_X4Y138_BO6),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_BLUT (
.I0(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_BQ),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_BQ),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.I4(CLBLL_L_X4Y137_SLICE_X4Y137_C5Q),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_DQ),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_ALUT (
.I0(CLBLM_R_X3Y138_SLICE_X3Y138_B5Q),
.I1(CLBLL_L_X2Y139_SLICE_X0Y139_BQ),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_B5Q),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_CQ),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_BO5),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_AO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_BO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_CO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_DLUT (
.I0(CLBLL_L_X2Y138_SLICE_X1Y138_AQ),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y138_SLICE_X1Y138_BQ),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccff00aaaa)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_CLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I1(CLBLM_R_X3Y138_SLICE_X3Y138_B5Q),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_B5Q),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccff00)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_BLUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ffcc00cc)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_AO5),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_CO5),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_AO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_CO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaa0a0a)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_DLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_CO6),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_A5Q),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_DO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccffcc00)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_CO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h888b888b88888888)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_BLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_BO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000ffaaaaf0f0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_B5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_AO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_CO5),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_DO5),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_AO6),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_BO6),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_CO6),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_DO6),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaffcc00ccff)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_DLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_DO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccffcc00)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_CLUT (
.I0(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_CQ),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y139_SLICE_X0Y139_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_CO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e0e0eeee)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_CQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_BO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00006a006a00)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I2(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_AO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_AO6),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_BO6),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_CO6),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_DO6),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0b1b1f5a0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I3(CLBLM_R_X3Y138_SLICE_X2Y138_CQ),
.I4(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I5(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f60606f505f505)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_CLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_C5Q),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ddf0ccf0ddf0cc)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_C5Q),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff0cccc00f0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_AO5),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_BO5),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_BO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_CO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_DO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000cffffaaaa)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_DLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_DO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_DO6),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0f0f0bbbb)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_CLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_CO6),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_CQ),
.I2(CLBLM_R_X7Y140_SLICE_X8Y140_B5Q),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505fa0acfc0cfc0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_BLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_CQ),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0f5fa050a)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_ALUT (
.I0(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.I1(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I4(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_AO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_BO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_CO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffffaf0f)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_DLUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_DQ),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_DQ),
.I3(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0aaf0aa)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_CLUT (
.I0(CLBLL_L_X4Y138_SLICE_X4Y138_AO6),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00008aba8aba)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_BLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_DQ),
.I1(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I2(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbf5515aaba0010)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I2(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I3(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I5(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X5Y141_AO6),
.Q(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500000005)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_DLUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_D5Q),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y61_I),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_C5Q),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc55dd00cc55dd)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_CLUT (
.I0(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.I1(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I4(CLBLM_R_X3Y139_SLICE_X3Y139_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000004055)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_CO6),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I3(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.I4(CLBLL_L_X4Y141_SLICE_X5Y141_CO6),
.I5(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fcfcfcfc)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I2(CLBLM_R_X5Y139_SLICE_X7Y139_DO6),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_C5Q),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_CO5),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_AO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a000a0000000000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_DLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y139_SLICE_X3Y139_C5Q),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555b88b8888)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_CLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf3fcfff0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_BLUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_CQ),
.I1(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_B5Q),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.I4(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc5acc5acc00cc00)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_ALUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_DO6),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_AO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_BO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffcc)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_C5Q),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I2(CLBLM_R_X3Y139_SLICE_X3Y139_C5Q),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I4(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3300aaaacc00)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_CO6),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b88bb888888888)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I4(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.I5(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_BO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1c0c0c00000ffff)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I3(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdccc100000550055)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_BLUT (
.I0(CLBLL_L_X4Y141_SLICE_X5Y141_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff5400fc0054)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I5(CLBLL_L_X4Y141_SLICE_X4Y141_CQ),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff0fff0fff)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fffffffc0000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_DO6),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc55ff550055)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_BLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_CQ),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3c00f000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_ALUT (
.I0(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_DO6),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_BO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_CO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_DO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fafaff003232)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_DLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe4fff000e400f0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_CLUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I5(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeefafa44445050)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbfaba55115010)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_CO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030fc30fc30)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf80d08fdf80d08)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_CLUT (
.I0(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaff88cc)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaafaf55000505)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_A5Q),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0101000051015000)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_B5Q),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afaff000ff0f)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_CLUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I4(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeaefea45404540)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I2(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_D5Q),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050dd88dd88)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_C5Q),
.I4(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_AO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_BO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffaaff30ffba)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_B5Q),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_DO6),
.I4(CLBLM_L_X8Y133_SLICE_X10Y133_CO6),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffffffefffff)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccccaaaa)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fafa5050)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0000000a880088)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_DLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_C5Q),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_BO6),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0c0cffff0c5d)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_CLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_C5Q),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_CO6),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_DO6),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbffff)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I3(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafc30ff00)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_AO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfcccfceefeeefe)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_CO6),
.I2(CLBLM_R_X3Y133_SLICE_X2Y133_B5Q),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_CO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y133_SLICE_X10Y133_BO6),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffbf)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_CLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7ffffffffbf)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaf0ccccaaaa)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_DQ),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeeefeeffffefee)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_DLUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_BO6),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcf00ccafefaaee)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_BO6),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaeaeffffffae)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_BLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_CO6),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_CO6),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_B5Q),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_DO6),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffffbff)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_ALUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_AO5),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_BO5),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_AO6),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_BO6),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00afaa0f00afaa)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_DLUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q),
.I4(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h083b000008080000)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_CLUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I4(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5a005accf0ccf0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_B5Q),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y134_SLICE_X13Y134_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3acacfc0cfc0c)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_DQ),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_AO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_BO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa0c0c0c0c)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_DLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.I3(1'b1),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0f4f0044)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_BO6),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.I4(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.I5(CLBLM_R_X7Y132_SLICE_X9Y132_CO6),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccccff00)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_BLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_DQ),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc55ccf0cc50)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_A5Q),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_AO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3fff33ff0fff00)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_CO6),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_BO5),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_B5Q),
.I5(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0000000a00)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_CLUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0022000000320010)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_CQ),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5a0f5a0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeeffffffcc)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_DO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_BO6),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff4444ffff44f4)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_CLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_D5Q),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.I4(CLBLM_L_X8Y135_SLICE_X11Y135_BO6),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000ba10)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I3(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffccceceffce)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_ALUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_BO6),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30baffff30ba30ba)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_DLUT (
.I0(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_CO6),
.I5(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeaffee)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_CLUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_BO6),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I2(CLBLM_L_X8Y132_SLICE_X10Y132_DO6),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_DO6),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_DO6),
.I5(CLBLM_L_X8Y136_SLICE_X10Y136_DO6),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000101010000000)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000000)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_ALUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_DQ),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_DO5),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_DO5),
.I4(CLBLM_L_X8Y137_SLICE_X10Y137_DO6),
.I5(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X11Y136_AO6),
.Q(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X11Y136_BO6),
.Q(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fafcfef0fafcfe)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_DLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_DQ),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_CO6),
.I4(CLBLM_L_X8Y138_SLICE_X11Y138_BO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff8a)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_CLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_DO6),
.I2(CLBLM_L_X10Y138_SLICE_X13Y138_AO6),
.I3(CLBLM_R_X7Y138_SLICE_X8Y138_CO6),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_DO6),
.I5(CLBLM_R_X7Y135_SLICE_X8Y135_CO6),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaf0f0cccc)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_BLUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfa00fafa)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_ALUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_D5Q),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_AO6),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000202000002020)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_DLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_DQ),
.I3(1'b1),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_DO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4040440040404400)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_CLUT (
.I0(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_CO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbaffbaffffffba)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_BLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I3(CLBLM_R_X7Y137_SLICE_X9Y137_BO6),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I5(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_BO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefaee50445044)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.I2(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_AO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_AO6),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_BO6),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00aaffffccee)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_DLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_CO6),
.I4(CLBLM_L_X8Y137_SLICE_X10Y137_CO6),
.I5(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_DO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h75ff757530ff3030)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_CLUT (
.I0(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_AO6),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_B5Q),
.I3(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_D5Q),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54aa00fe54fe54)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I2(CLBLM_L_X8Y134_SLICE_X10Y134_B5Q),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I5(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_BO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heceeeeec20222220)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_C5Q),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_AO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_B5Q),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300bbaabbaa)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_DLUT (
.I0(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.I2(1'b1),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_DO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8fff8fff8f8f8f8)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_CLUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_DO6),
.I3(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_CQ),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_CO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff303030)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y138_SLICE_X11Y138_BO6),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I5(CLBLM_R_X7Y138_SLICE_X8Y138_DO6),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_BO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbabaffba)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_DO6),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_CO6),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_AO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X11Y138_AO6),
.Q(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000585800000808)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_DLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_C5Q),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_DO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222f2f2ff22fff2)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_CLUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.I2(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_C5Q),
.I4(CLBLM_L_X8Y138_SLICE_X11Y138_BO5),
.I5(CLBLM_L_X12Y137_SLICE_X16Y137_AO6),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_CO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfffbfffffff)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_BO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fcfc5454)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_AQ),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_AO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_BO5),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_CO5),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_AO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_CO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8020080240100401)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_DLUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_C5Q),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ccccff00)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_CLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_C5Q),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00b1e4b1e4)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff0cccc5550)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_C5Q),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_CO5),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_DO5),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_AO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_BO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccff00)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccffcc00)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_C5Q),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaccaaf0aacc)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe3232ccfe0032)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I4(CLBLM_L_X8Y134_SLICE_X10Y134_B5Q),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_BO5),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_DO5),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_AO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_BO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_CO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_DO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0ee22ee22)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_DQ),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dd88dd88)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccffaaf0aaf0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_BLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I1(CLBLM_R_X3Y134_SLICE_X2Y134_DQ),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaffaac0aaf0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I5(CLBLM_R_X7Y140_SLICE_X8Y140_DQ),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_CO5),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_AO6),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_CO6),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_DO6),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf022f022f000f000)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_BO6),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccccf0ccf0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_CLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_D5Q),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_BQ),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccfff000cc00f0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ff55ea40fa50)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I5(CLBLM_R_X5Y139_SLICE_X6Y139_A5Q),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_BO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000011)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_DLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y138_SLICE_X7Y138_A5Q),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00fe54fe54)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7755070577550705)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_BO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa33aaf0aa30)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_ALUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_A5Q),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_DQ),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_AO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_B5Q),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_A5Q),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I4(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I5(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_BLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_AO5),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc5accffccf0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I5(CLBLM_L_X8Y141_SLICE_X11Y141_CO6),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f022222222)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000beeebeee)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_BLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_AO6),
.I4(CLBLL_L_X2Y137_SLICE_X0Y137_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heffeeffe23322332)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_ALUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_AO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050000050500000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I1(1'b1),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_ALUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_A5Q),
.I1(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0bff0fff04000000)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_DLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I5(CLBLM_R_X5Y143_SLICE_X7Y143_C5Q),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f373f37ff77ff77)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaccaaaa)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I2(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I3(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff70ff3400700034)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_DQ),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbf0000bfbf0000)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf020fffff000ffff)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0301ffff0303ffff)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_DQ),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_CO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_DO6),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ccccaaaa)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_CLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb51ab01fe54ae04)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I3(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_C5Q),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_DO6),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac0ccaaaaccc0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_ALUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_A5Q),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_A5Q),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb8b888bbbb888b8)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_ALUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I4(CLBLM_L_X10Y134_SLICE_X13Y134_CQ),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_CO6),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_DLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_CLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0070003000500000)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_BLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I5(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaff5000fa0050)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_A5Q),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_DLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080808088888888)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb0bfe0ef101f404)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_BLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y138_SLICE_X7Y138_A5Q),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_A5Q),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbb8b888bb88b8)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I3(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_AO5),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a2a200008080)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_B5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_B5Q),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_CLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_BO6),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_CO6),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_DO6),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_DO6),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff0200)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0aaf0aa)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_ALUT (
.I0(CLBLM_L_X10Y134_SLICE_X12Y134_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffeeee)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_DLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000000)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_DO6),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff0033ccfc0030)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_C5Q),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_BO5),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_AO6),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_BO6),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h11f1000000f00000)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_DLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I4(CLBLM_L_X12Y138_SLICE_X16Y138_AO6),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0105000501010000)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I4(CLBLM_L_X10Y137_SLICE_X12Y137_A5Q),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f055cc55cc55)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_BLUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaf05ccccfa50)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_CO5),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_AO6),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_BO6),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_CO6),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff02ff33ff02ff02)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_DLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_DO6),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccffcc00)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_CQ),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_A5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafc00fcfc)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_BLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_BQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccf0ccf0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I2(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I5(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_CO5),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_BO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_CO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddd8ddd888d888)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_DQ),
.I3(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30b8b8b8b8)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fe54ee44ae04)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_A5Q),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_A5Q),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fc000000fc)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.Q(CLBLM_L_X10Y135_SLICE_X13Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.Q(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.Q(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.Q(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff7f5f3f0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.I2(CLBLM_L_X10Y134_SLICE_X13Y134_DO6),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_DQ),
.I5(CLBLM_L_X8Y134_SLICE_X10Y134_CO6),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff31002000)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_R_X7Y137_SLICE_X9Y137_A5Q),
.I5(CLBLM_L_X10Y134_SLICE_X12Y134_CO6),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff000fc0cfc0cf)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I4(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cc0cfc0cf)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y137_SLICE_X9Y137_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_AO5),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_AO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_BO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000083838080)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_B5Q),
.I5(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfffffffffbffff)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaff3c003c)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_BLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_CQ),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y139_SLICE_X13Y139_DQ),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc303088bb88bb)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_ALUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_CO6),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.Q(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0031ffff0031)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_DLUT (
.I0(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_DO6),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.I3(CLBLM_R_X11Y136_SLICE_X14Y136_AO5),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f400f700f000f0)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_CLUT (
.I0(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_BO6),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_CO6),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I5(CLBLM_L_X12Y137_SLICE_X16Y137_CO6),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000c00080000)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbbfbffffaafa)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_ALUT (
.I0(CLBLM_L_X10Y137_SLICE_X13Y137_DO6),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_D5Q),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_AO6),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_CO6),
.I5(CLBLM_R_X3Y137_SLICE_X2Y137_CQ),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_AO6),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696696969699696)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.I1(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I2(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I5(CLBLM_L_X10Y137_SLICE_X12Y137_BO6),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffffffffffe)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55acc00ff33)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_BLUT (
.I0(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ffcc00ccff)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_C5Q),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff4fff444444444)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h02028a0200008800)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_CQ),
.I4(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.I5(CLBLM_L_X10Y134_SLICE_X13Y134_C5Q),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff7530)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_BLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_CO6),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_AO6),
.I2(CLBLM_L_X10Y134_SLICE_X13Y134_C5Q),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_CQ),
.I4(CLBLM_L_X10Y137_SLICE_X13Y137_AO6),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_DO6),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d0c5d0cffff5d0c)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_ALUT (
.I0(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_A5Q),
.I4(CLBLM_L_X10Y137_SLICE_X13Y137_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_BO6),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_CO6),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_DO6),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888d8d8d8d8)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I5(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f0fcccc00ff)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_CLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I1(CLBLM_R_X3Y138_SLICE_X2Y138_BQ),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0aaaaff00)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_BLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.I1(1'b1),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3f3aaaac0c0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.Q(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff75ff30)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_DLUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I5(CLBLM_L_X10Y138_SLICE_X13Y138_BO6),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffbf0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_CLUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_AO6),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_DO6),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_DO6),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I4(CLBLM_L_X10Y138_SLICE_X13Y138_DO6),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_DO6),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000800)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_C5Q),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0500ffff1100)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_ALUT (
.I0(CLBLM_R_X11Y138_SLICE_X14Y138_DO6),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.I2(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I3(CLBLM_R_X11Y138_SLICE_X14Y138_BO6),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_BO6),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y137_SLICE_X2Y137_CQ),
.Q(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_CQ),
.Q(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5dff0cff5d5d0c0c)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_A5Q),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_AO6),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_CO6),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_DO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7fffffffff7)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffffffcfc)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_BLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_DQ),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_BO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcf030300aa0055)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_ALUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_AO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_AO5),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X14Y139_CO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_CO5),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_AO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_BO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_CO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_DO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0a0f5b1a0e4f5)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.I4(CLBLM_L_X10Y137_SLICE_X12Y137_DO6),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_DO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0d8d8d8d8)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_C5Q),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_CO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe0e0ef0fe000e)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_DQ),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_CQ),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_BO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfafa0a0a)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_ALUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_CO6),
.I1(CLBLM_R_X11Y137_SLICE_X15Y137_AO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I4(CLBLM_R_X3Y133_SLICE_X2Y133_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_AO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_AO5),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_AO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X14Y140_AO5),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_AO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_BO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_CO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h09cc0ccc55005500)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_DLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_DO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefab4501feba5410)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.I3(CLBLM_L_X8Y140_SLICE_X11Y140_C5Q),
.I4(CLBLM_R_X5Y140_SLICE_X7Y140_B5Q),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_CO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fefc0e0c)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_BLUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.I4(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_BO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_ALUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_BO6),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_AO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_C5Q),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_DO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff7fffffff)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_CO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7070705200220022)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_BLUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_BO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0d1e2aa00aa00)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_ALUT (
.I0(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_B5Q),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_AO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_AO6),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_BO6),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080000000000000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_DLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AO5),
.I3(1'b1),
.I4(CLBLM_L_X10Y141_SLICE_X12Y141_BQ),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_AO6),
.I4(CLBLM_L_X10Y141_SLICE_X12Y141_DO6),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ae04ff55ff55)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_BQ),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_C5Q),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_CO6),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc50cc50cc50)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_ALUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_AO5),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_CO5),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_AO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_BO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_DLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_C5Q),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ccccaa00aaf0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_CLUT (
.I0(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I1(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y141_SLICE_X11Y141_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b8b888b88888b88)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_BLUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.I4(CLBLM_L_X8Y141_SLICE_X11Y141_BO6),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000007878)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_ALUT (
.I0(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_B5Q),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I3(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_BO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080000080800000)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_AO6),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf3aaf3aafcaafc)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd8dd88833333333)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I3(CLBLM_R_X11Y141_SLICE_X14Y141_CO6),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000000000000)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_DLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_C5Q),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1555555555555555)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_CLUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_AO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_C5Q),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_DO5),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffec00ecff200020)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_BLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_DO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_A5Q),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_CO6),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa00faff0a000a)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y134_SLICE_X13Y134_C5Q),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_CO6),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.Q(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.Q(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_CO6),
.Q(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0fc00cc)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccffa000a0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_BLUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_DO6),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_CO6),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y140_SLICE_X7Y140_C5Q),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccf0ccaaccaa)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_CO5),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_AO6),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_BO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h07770fff0fff0fff)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_DLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I4(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff7fffffff)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffcc00aa00cc)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_C5Q),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa000a0ffac00ac)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_DO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_A5Q),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_ALUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff7fffff)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_BLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffeffffffffff)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_ALUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_DO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_CO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefffff)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_BO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff0000a088)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_DO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_CO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_BO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_AO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0f0f0)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_DLUT (
.I0(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_BO6),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_DO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000080c00000a0f0)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_CLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_BO6),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_CO6),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_DQ),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_BO5),
.I5(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_CO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffeeff00310020)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_BO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdffffffffffff7)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_DO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_CO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_BO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcccf000fcccf000)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_AO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heca0eca0eca0eca0)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_DLUT (
.I0(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_CQ),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_DO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000d0dd)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X11Y138_SLICE_X14Y138_AO5),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.I3(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I4(CLBLM_L_X12Y138_SLICE_X16Y138_BO5),
.I5(CLBLM_R_X11Y139_SLICE_X14Y139_DO5),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_CO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ffff00200000)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_BO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005522200020)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I2(RIOB33_X105Y137_IOB_X1Y138_I),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_R_X7Y139_SLICE_X8Y139_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_AO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_DO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_CO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_BO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_AO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_DO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_CO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_BO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333bbbbbbbb)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X13Y138_CO6),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y135_SLICE_X14Y135_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_AO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_DO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_CO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_BO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33ff33ff33)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_AO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X3Y129_BO6),
.Q(CLBLM_R_X3Y129_SLICE_X3Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X3Y129_AO6),
.Q(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aac0c00000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_BLUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaafaa05000500)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y138_SLICE_X2Y138_CQ),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000088008800)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000cccc0000cccc)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_ALUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_A5Q),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffcc)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y134_SLICE_X3Y134_CQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y132_SLICE_X3Y132_A5Q),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I5(CLBLM_R_X3Y133_SLICE_X2Y133_BQ),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff00ff01)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_CLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_B5Q),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_D5Q),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_DO6),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc5554fffc5555)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_BLUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_BO5),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_BO6),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_A5Q),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_D5Q),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_CO6),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5f0f0fff5fcf4)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_DO6),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_D5Q),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_C5Q),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_CO6),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_AO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3a0a0fa0afa0a)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_ALUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_AO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_AO5),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_AO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ff66ff66ff66ff6)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_DLUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_A5Q),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I2(CLBLM_R_X3Y133_SLICE_X2Y133_B5Q),
.I3(CLBLM_R_X3Y132_SLICE_X3Y132_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00408840)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_CLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_D5Q),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_A5Q),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_DO6),
.I5(CLBLM_R_X3Y132_SLICE_X3Y132_BO6),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h001b0000000a0000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_BLUT (
.I0(CLBLM_R_X3Y140_SLICE_X3Y140_A5Q),
.I1(CLBLL_L_X4Y137_SLICE_X4Y137_D5Q),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0aaccaacc)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_ALUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_B5Q),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X2Y133_BO5),
.Q(CLBLM_R_X3Y133_SLICE_X2Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X2Y133_CO5),
.Q(CLBLM_R_X3Y133_SLICE_X2Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X2Y133_AO6),
.Q(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X2Y133_BO6),
.Q(CLBLM_R_X3Y133_SLICE_X2Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X2Y133_CO6),
.Q(CLBLM_R_X3Y133_SLICE_X2Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2020a000a0a00000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_DLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_DO6),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ffaa5500)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I2(LIOB33_X0Y63_IOB_X0Y63_I),
.I3(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacfc0cfc0c)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_BLUT (
.I0(CLBLL_L_X2Y139_SLICE_X1Y139_CQ),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdd00ddffd000d0)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_C5Q),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_BO5),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_A5Q),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_BO6),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ccf5ccf5)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_CLUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_C5Q),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I2(CLBLM_R_X3Y133_SLICE_X2Y133_DO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_BO6),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f055ff550055)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_BLUT (
.I0(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I1(1'b1),
.I2(CLBLM_R_X3Y139_SLICE_X3Y139_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc50cc00cc00cc00)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_ALUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X3Y140_A5Q),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X2Y135_AO6),
.Q(CLBLM_R_X3Y134_SLICE_X2Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X2Y134_AO6),
.Q(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X2Y134_BO6),
.Q(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X2Y134_CO6),
.Q(CLBLM_R_X3Y134_SLICE_X2Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X2Y134_DO6),
.Q(CLBLM_R_X3Y134_SLICE_X2Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d8d8d8d8)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_DLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I1(CLBLM_R_X3Y134_SLICE_X2Y134_CQ),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_DO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa800a8fffc00fc)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_CLUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I1(CLBLM_R_X3Y134_SLICE_X2Y134_CQ),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.I5(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_CO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000006c006c)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_BLUT (
.I0(CLBLM_R_X3Y135_SLICE_X2Y135_CO6),
.I1(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_DQ),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_BO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000012121212)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_ALUT (
.I0(CLBLM_R_X3Y135_SLICE_X2Y135_CO6),
.I1(CLBLM_R_X3Y134_SLICE_X3Y134_DQ),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_AO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_CO5),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_DO5),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_AO6),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_BO6),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_CO6),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_DO6),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0fcfc0c0c)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_DLUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_A5Q),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_DO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0dddd8888)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_D5Q),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_B5Q),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_CO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f9f9f9f9)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_CO6),
.I1(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I3(CLBLM_R_X3Y134_SLICE_X2Y134_A5Q),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_BO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888b888b88b888b8)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_DQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y135_SLICE_X2Y135_AO5),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_AO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.Q(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.Q(CLBLM_R_X3Y135_SLICE_X2Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_DO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_CLUT (
.I0(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_BQ),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I3(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I5(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_CO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h888800007fff7fff)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_BLUT (
.I0(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I1(CLBLM_R_X3Y134_SLICE_X2Y134_BQ),
.I2(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I3(CLBLL_L_X2Y135_SLICE_X1Y135_DQ),
.I4(CLBLM_R_X3Y135_SLICE_X2Y135_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_BO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888a000a000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I4(CLBLL_L_X2Y139_SLICE_X0Y139_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_AO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_CO5),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_AO6),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_BO6),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_CO6),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_DO6),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hababbaba01011010)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y134_SLICE_X3Y134_DQ),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I5(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_DO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ccccff00)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_CLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I1(CLBLM_R_X3Y134_SLICE_X2Y134_CQ),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_A5Q),
.I3(CLBLL_L_X4Y135_SLICE_X5Y135_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_CO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ccccf000)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I3(CLBLL_L_X2Y135_SLICE_X1Y135_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X2Y135_SLICE_X1Y135_BQ),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_BO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffaf00ef00af)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.I1(CLBLL_L_X2Y135_SLICE_X1Y135_AQ),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y135_SLICE_X1Y135_BQ),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_AO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_AO6),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_BO6),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_CO6),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000005fffffff)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_DLUT (
.I0(CLBLM_R_X3Y136_SLICE_X2Y136_BQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I4(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_DO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000012221222)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_CLUT (
.I0(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I1(CLBLM_R_X3Y134_SLICE_X3Y134_DQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I4(CLBLM_R_X3Y137_SLICE_X2Y137_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_CO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a3acacac)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_BLUT (
.I0(CLBLM_R_X3Y138_SLICE_X3Y138_DQ),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I4(CLBLM_R_X3Y135_SLICE_X2Y135_AO5),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_DQ),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_BO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddccdd00110011)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_ALUT (
.I0(CLBLM_R_X3Y135_SLICE_X2Y135_BO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y136_SLICE_X2Y136_DO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_BQ),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_AO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_AO5),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_BO5),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_CO5),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_DO5),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_AO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_BO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_CO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_DO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f20202fc0cfc0c)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_DLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.I4(CLBLM_R_X3Y133_SLICE_X2Y133_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_DO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c5c5f505f505)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X2Y139_SLICE_X1Y139_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_CO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccf0ccf0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_BO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccfff000f0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_ALUT (
.I0(CLBLM_R_X3Y140_SLICE_X3Y140_C5Q),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_AO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X2Y137_DO5),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X2Y137_AO6),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X2Y137_BO6),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X2Y137_CO6),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X2Y137_DO6),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2dd11dd11)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_DLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I3(CLBLM_R_X3Y138_SLICE_X2Y138_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_DO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55af05ee44ae04)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y137_SLICE_X2Y137_CQ),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I3(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I5(CLBLL_L_X4Y135_SLICE_X5Y135_A5Q),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_CO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccac0000ccac)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_BLUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I1(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.I2(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I3(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y137_SLICE_X3Y137_B5Q),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_BO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333dffd1331)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_ALUT (
.I0(CLBLM_R_X3Y135_SLICE_X2Y135_BO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I3(CLBLM_R_X3Y136_SLICE_X2Y136_DO6),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_CQ),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_DQ),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_AO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_BO5),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_CO5),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_DO5),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_AO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_BO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_CO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_DO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3c0b8b8b8b8)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_DLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X2Y137_SLICE_X1Y137_C5Q),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_C5Q),
.I4(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_DO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaafff000f0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_CLUT (
.I0(LIOB33_X0Y59_IOB_X0Y59_I),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_CO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fc0cfc0c)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_DQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_B5Q),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_BO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffd000dd00d0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y134_SLICE_X3Y134_D5Q),
.I5(CLBLL_L_X2Y139_SLICE_X1Y139_DQ),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_AO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X2Y138_AO5),
.Q(CLBLM_R_X3Y138_SLICE_X2Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X2Y138_AO6),
.Q(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X2Y138_BO6),
.Q(CLBLM_R_X3Y138_SLICE_X2Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X2Y138_CO6),
.Q(CLBLM_R_X3Y138_SLICE_X2Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X2Y138_DO6),
.Q(CLBLM_R_X3Y138_SLICE_X2Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3cff3c003c003c)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y59_IOB_X0Y60_I),
.I2(CLBLM_R_X3Y138_SLICE_X2Y138_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_DO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ddf0fff000f022)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_CLUT (
.I0(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I1(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I5(CLBLM_R_X3Y137_SLICE_X2Y137_BQ),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_CO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffafffaf)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_BLUT (
.I0(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I2(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_BO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa0fffaa00aa)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_ALUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_AO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_AO5),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_BO5),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_CO5),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_DO5),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_AO6),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_BO6),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_CO6),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_DO6),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333aaaa3333)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_DLUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y137_SLICE_X4Y137_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_DO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcffc0330bbbb8888)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_CLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_D5Q),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I4(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_CO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f606fff00f00)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_BLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X2Y139_SLICE_X0Y139_BQ),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_BO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88cffc0330)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_ALUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_AO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y140_SLICE_X2Y140_BQ),
.Q(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h333300000f000f00)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_B5Q),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I4(CLBLM_R_X3Y139_SLICE_X3Y139_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_DO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44440000c0c00000)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_CLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I2(CLBLL_L_X2Y139_SLICE_X1Y139_BQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y139_SLICE_X1Y139_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_CO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fffffff7ffffff)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_BLUT (
.I0(CLBLL_L_X2Y139_SLICE_X1Y139_BQ),
.I1(CLBLL_L_X2Y139_SLICE_X1Y139_CQ),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I3(CLBLL_L_X2Y139_SLICE_X1Y139_DQ),
.I4(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd8d8800ffff00)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y139_SLICE_X3Y139_B5Q),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_BQ),
.I3(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I4(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X2Y139_AO6),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X3Y139_BO5),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X3Y139_CO5),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X3Y139_AO6),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X3Y139_BO6),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X3Y139_CO6),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5855505555555555)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_DLUT (
.I0(CLBLM_R_X3Y139_SLICE_X3Y139_C5Q),
.I1(CLBLL_L_X2Y139_SLICE_X1Y139_DQ),
.I2(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I4(CLBLM_R_X3Y139_SLICE_X2Y139_CO5),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_DO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee228888b8b8)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_CLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I4(CLBLM_R_X3Y139_SLICE_X3Y139_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_CO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00e4e4e4e4)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y138_SLICE_X3Y138_DQ),
.I2(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_BO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff55ccccf050)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I1(CLBLM_R_X3Y139_SLICE_X3Y139_BQ),
.I2(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y138_SLICE_X2Y138_A5Q),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_AO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X2Y140_CO6),
.Q(CLBLM_R_X3Y140_SLICE_X2Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X2Y140_AO6),
.Q(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X2Y140_BO6),
.Q(CLBLM_R_X3Y140_SLICE_X2Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a0a0a0a0a)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_DO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff33ff33ff33)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_CLUT (
.I0(CLBLM_R_X3Y138_SLICE_X3Y138_A5Q),
.I1(CLBLM_R_X3Y139_SLICE_X3Y139_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X3Y135_SLICE_X2Y135_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_CO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffaaba45550010)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I2(CLBLL_L_X2Y137_SLICE_X1Y137_BQ),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I5(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_BO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd88dd88d88888888)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_AO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_AO5),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_CO5),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_AO6),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_BO6),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_CO6),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ffffffa0000000)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_DO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3acacfa0afa0a)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_CLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_C5Q),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_B5Q),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_DO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_CO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd9ff9900d90099)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_BLUT (
.I0(CLBLM_R_X3Y140_SLICE_X3Y140_DO6),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.I2(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(LIOB33_X0Y55_IOB_X0Y55_I),
.I5(CLBLM_R_X3Y138_SLICE_X3Y138_CQ),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_BO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffaa00aa)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_ALUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_CO6),
.I1(CLBLM_R_X3Y141_SLICE_X3Y141_CO6),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_AO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.Q(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.Q(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff101400001014)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_B5Q),
.I1(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_DQ),
.I3(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfaafccccfafa)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_ALUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_B5Q),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y141_SLICE_X2Y141_CO6),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y141_SLICE_X3Y141_AO6),
.Q(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y141_SLICE_X3Y141_BO6),
.Q(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccccccccccc)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.I1(LIOB33_X0Y55_IOB_X0Y55_I),
.I2(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_C5Q),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.I5(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf3fc0c03f3fc0c0)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_CLUT (
.I0(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_C5Q),
.I3(LIOB33_X0Y55_IOB_X0Y55_I),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0b1e4a0a0a0e4)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_BQ),
.I3(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_B5Q),
.I5(CLBLL_L_X4Y141_SLICE_X4Y141_DQ),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dd888888dd88888)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.I2(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.Q(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50fe54ba10)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y165_SLICE_X2Y165_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y165_SLICE_X2Y165_DO5),
.O6(CLBLM_R_X3Y165_SLICE_X2Y165_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y165_SLICE_X2Y165_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y165_SLICE_X2Y165_CO5),
.O6(CLBLM_R_X3Y165_SLICE_X2Y165_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y165_SLICE_X2Y165_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y165_SLICE_X2Y165_BO5),
.O6(CLBLM_R_X3Y165_SLICE_X2Y165_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_R_X3Y165_SLICE_X2Y165_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y165_SLICE_X2Y165_AO5),
.O6(CLBLM_R_X3Y165_SLICE_X2Y165_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y165_SLICE_X3Y165_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y165_SLICE_X3Y165_DO5),
.O6(CLBLM_R_X3Y165_SLICE_X3Y165_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y165_SLICE_X3Y165_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y165_SLICE_X3Y165_CO5),
.O6(CLBLM_R_X3Y165_SLICE_X3Y165_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y165_SLICE_X3Y165_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y165_SLICE_X3Y165_BO5),
.O6(CLBLM_R_X3Y165_SLICE_X3Y165_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y165_SLICE_X3Y165_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y165_SLICE_X3Y165_AO5),
.O6(CLBLM_R_X3Y165_SLICE_X3Y165_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_CO5),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_CLUT (
.I0(RIOB33_X105Y123_IOB_X1Y123_I),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I2(CLBLM_L_X8Y134_SLICE_X10Y134_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000a3aca3ac)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_BLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_DQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_DO6),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fafa5050)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c00000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c0c000000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_CO5),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_DO5),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_DO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc33008b8b8888)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_DLUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_D5Q),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaccfff000f0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_CLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00bebebebe)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_BLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffc000000fc)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_B5Q),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_CO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3fffffffffffff)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000f0f0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_DQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff66f0f0ff66)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aafcaaf0aa30)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_DO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_BO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0e2aa00aa00)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_DLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_B5Q),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff10ff4000100040)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_DO5),
.I5(CLBLM_R_X3Y135_SLICE_X2Y135_BQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f6fcf6fc)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_DO6),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbeafbea51405140)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y135_SLICE_X1Y135_CQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b7b7b7bdededede)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_DLUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_CQ),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_D5Q),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fbfdfef7fbfdfe)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_CLUT (
.I0(CLBLM_R_X3Y133_SLICE_X2Y133_BQ),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_C5Q),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_DO6),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbeffffbe)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_BLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_B5Q),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_CQ),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_B5Q),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc5acc00cc5a)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I5(CLBLL_L_X4Y136_SLICE_X4Y136_B5Q),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_AO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_BO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_CO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_DO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00d8d8d8d8)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_DLUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.I2(CLBLM_R_X5Y133_SLICE_X6Y133_DQ),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ff55ee44aa00)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I5(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacfcacacac0ca)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_BLUT (
.I0(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00c8c8fafa)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_ALUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_BO5),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_CO5),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_DO5),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_AO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_BO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb88bbc0f3c0f3)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222ee22ee22)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_CLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y133_SLICE_X2Y133_C5Q),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0f000ff0f)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_BLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_CQ),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0fff000f0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_CO5),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_BO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_CO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_DO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d888dddddd)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88ff33cc00)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y135_SLICE_X1Y135_DQ),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb88bbdede1212)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I4(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff003030)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_CO5),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_DO5),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_AO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_BO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_CO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11ee44e4e4e4e4)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_B5Q),
.I3(CLBLM_R_X3Y138_SLICE_X2Y138_DQ),
.I4(CLBLM_R_X7Y140_SLICE_X9Y140_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44afaf0505)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y133_SLICE_X2Y133_BQ),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f5c4f5c4)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_BLUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_D5Q),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccf5cc00cca0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I2(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I5(CLBLM_R_X5Y136_SLICE_X7Y136_A5Q),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_CO5),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_DO5),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_BO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_CO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_DO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0f3f3cd01cd01)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_DLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y135_SLICE_X4Y135_CQ),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y135_SLICE_X5Y135_A5Q),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeff0e0ff2f00200)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_BLUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.I5(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff600f6ff000000)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_C5Q),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y135_SLICE_X1Y135_BQ),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_A5Q),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ff66ff66ff66ff6)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_DLUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_A5Q),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000909000000909)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_CLUT (
.I0(CLBLM_R_X7Y140_SLICE_X9Y140_D5Q),
.I1(CLBLL_L_X2Y135_SLICE_X1Y135_DQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_DO6),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3acacff0ff000)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_A5Q),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_B5Q),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3333aaaa3030)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X6Y133_DQ),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_BO5),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_CO5),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_DO5),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_AO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_BO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_CO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_DO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaff00cccc)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_DLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccf0f0aaaa)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_CLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_D5Q),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_D5Q),
.I2(CLBLM_R_X3Y137_SLICE_X2Y137_BQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc55aaf0f0cccc)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_BLUT (
.I0(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_BQ),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafff0aaaa3330)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_D5Q),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_AO5),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_BO5),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_CO5),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_AO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_BO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_CO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaeeffff00cc)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_DLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_DO6),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1b1b1bb11bb11)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_C5Q),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000acacacac)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_BLUT (
.I0(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y141_SLICE_X12Y141_BQ),
.I4(RIOB33_X105Y123_IOB_X1Y124_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303fc0cacacacac)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I4(CLBLM_R_X5Y140_SLICE_X6Y140_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_BO5),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_CO5),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_BO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_CO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00dd88dd88)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5a5aff00aaaa)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_CQ),
.I2(CLBLL_L_X4Y135_SLICE_X4Y135_B5Q),
.I3(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_CO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dddd88e4e4e4e4)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_BO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fffa5550)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_DQ),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_AO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_CO5),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_AO6),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_BO6),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_CO6),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3020002030200020)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_DLUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_DO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaff00cccc)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_B5Q),
.I3(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_CO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfff00f00)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X2Y137_SLICE_X1Y137_AQ),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.I5(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_BO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3f3aaaaf300)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_ALUT (
.I0(CLBLM_R_X7Y140_SLICE_X9Y140_DQ),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_AO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_BO5),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_CO5),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_AO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_CO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffefffe)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_B5Q),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_CQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f3f3c0ee22ee22)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ccaaccaa)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_BLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_D5Q),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccfff000f0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_A5Q),
.I5(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_AO5),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_CO5),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_AO6),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_BO6),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_CO6),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050004400500044)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_DLUT (
.I0(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.I2(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbebe1414ee44ee44)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I2(CLBLL_L_X4Y135_SLICE_X4Y135_DQ),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bb88bb8eeee2222)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_BLUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_C5Q),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3acacfa0afa0a)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_ALUT (
.I0(CLBLM_R_X5Y138_SLICE_X7Y138_B5Q),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_DQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_AO5),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_AO6),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_CO6),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfc)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y138_SLICE_X3Y138_A5Q),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X5Y140_SLICE_X7Y140_CQ),
.I5(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888b8888888b)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_CLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3d1c0c0c0c0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_BLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I3(CLBLL_L_X4Y134_SLICE_X5Y134_CO6),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5050f0f0ff00)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_ALUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_DQ),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_A5Q),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_AO6),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_BO6),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_CO6),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffdfe)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_DLUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_BO6),
.I2(CLBLM_R_X7Y139_SLICE_X8Y139_DO6),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_DO6),
.I5(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d888d8d88dd8888)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_BO5),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_B5Q),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf5f0cccc5500)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_BLUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_BO5),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I2(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.I3(CLBLL_L_X4Y141_SLICE_X4Y141_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00acacacac)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_ALUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_AO5),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_BO5),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_CO5),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_BO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_CO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_BQ),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_A5Q),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_D5Q),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_DO6),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50b1b1b1b1)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_BQ),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0fafa0a0a)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_DQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I4(CLBLM_R_X5Y140_SLICE_X7Y140_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f03333ff00cccc)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_BO5),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_CO5),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_DO5),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_AO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_BO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_CO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_DO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_CQ),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0ff0ccccff00)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_CLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_C5Q),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.I2(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccccccaaaa)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00bbbbb0b0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_DQ),
.I4(CLBLM_R_X5Y140_SLICE_X7Y140_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_BO5),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_CO5),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_AO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_BO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_CO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h555541550000ff00)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_DLUT (
.I0(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_C5Q),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_C5Q),
.I3(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cafa0afa0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_CLUT (
.I0(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0ee22ee22)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y139_SLICE_X3Y139_C5Q),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I4(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd01dc10ef23fe32)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_DO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.I4(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I5(CLBLM_L_X10Y131_SLICE_X12Y131_C5Q),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.Q(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X7Y141_BO6),
.Q(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ff66ffff66ff66)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_DLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_DQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a000a000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I3(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aaccaacc)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_BLUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_DQ),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc50cca0cc50cca0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_CQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_AO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_BO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222222222222)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_DLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_C5Q),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4f5e4f5b1f5b1)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y134_SLICE_X5Y134_DO6),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff55cc44)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_BLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cc00fc30cc00)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I5(CLBLM_R_X5Y141_SLICE_X7Y141_CO6),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_DO5),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_AO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_BO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_DO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0acfcfc0c0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_DLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_D5Q),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4fa50fa50)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_D5Q),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_C5Q),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfc0d0cf8fc080c)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_C5Q),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ea40ff55fa50)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_C5Q),
.I5(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_DO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_BO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_CO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f70007)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_C5Q),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0ffe0efe0e)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_BLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0cfcfcfcf)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y134_SLICE_X5Y134_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_CO5),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff80008080808080)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y141_SLICE_X5Y141_DO6),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_A5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaccccf0f0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f022882288)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_BLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff002828ff00a0a0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_AO5),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_AO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22bbbb8888)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_ALUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccffcc00)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_D5Q),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I2(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000000f0f00000)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_DO6),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_CLUT (
.I0(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_DO6),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfeabae51540104)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_DO5),
.I4(CLBLM_R_X3Y134_SLICE_X3Y134_C5Q),
.I5(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdcdfece31013202)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_C5Q),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_B5Q),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_CO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ccffcc55)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0aaf0aa)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff3000330030)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X3Y140_A5Q),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_BO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_DO6),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00cfcfc0c0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I4(CLBLM_R_X3Y138_SLICE_X3Y138_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa3ffac00a300ac)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_A5Q),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_BQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00bebeff001414)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_C5Q),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_B5Q),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_DLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_BQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_CLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0ffaa5500)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I3(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22bbb88b88)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_ALUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_BO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000aa0c000c00)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_DLUT (
.I0(CLBLM_R_X3Y138_SLICE_X3Y138_C5Q),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000100022000000)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_CO6),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f3c0f3ccff0033)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeff4455eafa4050)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I4(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I5(CLBLL_L_X4Y133_SLICE_X5Y133_CQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa000020202020)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_DLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_BO6),
.I2(CLBLL_L_X4Y137_SLICE_X5Y137_CQ),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000500033000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_CO5),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_BO6),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_DQ),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_R_X3Y137_SLICE_X2Y137_DQ),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h220000002200a0a0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_CO5),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_A5Q),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_A5Q),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_BO6),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_DO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_BO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_CO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0c00008888)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_DLUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01100f0f04400)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_DO5),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aafff0f088cc)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_CQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_A5Q),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0fcc00ccf0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_D5Q),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_CO5),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_BO5),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002320)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_DLUT (
.I0(CLBLM_R_X3Y135_SLICE_X2Y135_BQ),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_DQ),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffeeffff0ff000)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I1(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000cfcfc0c0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_CQ),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd01ce02ce02ce02)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_C5Q),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_DO5),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_AO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_BO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_CO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_DO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ffaa5500)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_B5Q),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I4(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ff55ea40ee44)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_D5Q),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_D5Q),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccfff000f0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaff3200fa0032)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_ALUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_A5Q),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_BO5),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_DO5),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_AO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_BO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_CO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_DO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ccaaccaa)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_DLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_C5Q),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff230023)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I1(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_D5Q),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0cc5acc5a)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_BLUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000a8fca8fc)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I1(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000002c200000)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_DLUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I3(CLBLM_R_X5Y140_SLICE_X6Y140_C5Q),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_CO6),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaafaeefe)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_CLUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_DO6),
.I1(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_CO6),
.I4(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.I5(CLBLM_R_X7Y135_SLICE_X8Y135_BO6),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbfabbaabbaa)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_BLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_DO6),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_AO6),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_D5Q),
.I4(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000000000)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_ALUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_C5Q),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_AO5),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_AO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_BO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fff3f3f0fff0f0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_CO6),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_BO5),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_B5Q),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafefafafafa)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I2(CLBLM_L_X8Y130_SLICE_X11Y130_AO6),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_DQ),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000f0ccf000)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_CO6),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00aaffaa00)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_ALUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_AO5),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_BO5),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_AO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_BO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7373ffff5050)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_CO6),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_CO6),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_DQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000000)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_CLUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_BO6),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_AO6),
.I5(CLBLM_R_X7Y135_SLICE_X8Y135_AO6),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaaaccaacc)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_BLUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_D5Q),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e288bb8888)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_ALUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_CQ),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_CO5),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_AO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_BO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff3fffffff0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_DO6),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_DO6),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf0aaf0aa)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa00aafc)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_BLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22dd11de12)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_ALUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_BO5),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_CO5),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_AO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_BO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_CO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcccceeffeeee)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I5(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccff660066)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_CLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0fff000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_BLUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa5550bbba1110)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_AO5),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_AO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3fff3f0f0fff0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y137_SLICE_X16Y137_AO6),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_CO6),
.I5(CLBLM_R_X3Y137_SLICE_X2Y137_D5Q),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fcf0fcfafefafe)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_CLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_CO6),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_BO6),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000008)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_BLUT (
.I0(CLBLM_R_X7Y140_SLICE_X9Y140_DQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afcfc0c0c)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_B5Q),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_A5Q),
.I4(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_AO5),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_AO6),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_BO6),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000af000000a0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_C5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.I5(CLBLM_R_X3Y138_SLICE_X3Y138_D5Q),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_DO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faf0fafffff0fa)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_CLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_DO6),
.I3(CLBLM_L_X12Y137_SLICE_X16Y137_AO6),
.I4(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_CO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ffd800d8)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_BLUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_BO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ff005a5a)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_ALUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I3(CLBLM_R_X3Y138_SLICE_X3Y138_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_AO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_AO6),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ffff33ccffffcc)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_A5Q),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_DO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d5dff5d0c0cff0c)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_CLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_CO6),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_DQ),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_CO6),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.I5(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_CO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffc0cf000fc0c)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_BO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbffb000bb00b0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_CQ),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_AO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.Q(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.Q(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.Q(CLBLM_R_X7Y139_SLICE_X8Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff5affa5ff5affa)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_DLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080808000000000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_CLUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_AO6),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff6ff6ffff6ff6)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_C5Q),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I4(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.I4(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X12Y139_AO6),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_AO6),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77dd77ddbbeebbee)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfffffffeff)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_CLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_DO6),
.I2(CLBLL_L_X4Y135_SLICE_X5Y135_DO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_DO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I5(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccec00000020)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_DQ),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfc0cfcfc0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q),
.I4(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_CO6),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_BO5),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_DO5),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_AO6),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_BO6),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_CO6),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_DO6),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0bbee1144)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_B5Q),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aaccaacc)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_CLUT (
.I0(CLBLM_R_X7Y137_SLICE_X8Y137_C5Q),
.I1(CLBLM_R_X7Y140_SLICE_X8Y140_CQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000acacacac)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_BLUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_CQ),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfaccfacc00ccfa)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_ALUT (
.I0(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_C5Q),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_CO5),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_DO5),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_AO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_BO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_CO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cfc0cfc0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_DLUT (
.I0(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44eeee4444)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X8Y140_SLICE_X11Y140_DQ),
.I4(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fcaaaa00fc)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_BLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I3(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccccf0cc)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.I2(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X8Y141_DO5),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X8Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X8Y141_BO6),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X8Y141_CO6),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0decc1200)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_DLUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_AO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I4(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffebee0000ebee)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_D5Q),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_CQ),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_DO6),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff006060c0c0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_BLUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_A5Q),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caaf0aa00aa00)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_ALUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_CO5),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_CO5),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_DO5),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_BO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_CO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_DO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ffcc00cc)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_DLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300e2e2e2e2)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_CLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y140_SLICE_X8Y140_DQ),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff1100ff0011)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_B5Q),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000078007800)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_ALUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_AO6),
.I2(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I4(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_CO5),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001110000)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_A5Q),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X4Y141_SLICE_X5Y141_DO6),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_B5Q),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X3Y139_SLICE_X3Y139_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8fa080afaf80a08)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_BLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_A5Q),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_D5Q),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3a3a3f303f303)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_ALUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_CQ),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff6cffccffccffcc)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_DLUT (
.I0(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_A5Q),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_B5Q),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_B5Q),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0a0000003133)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_DQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I3(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaa3300)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_B5Q),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ff00b8b8)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_CO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00020230303030)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y141_SLICE_X5Y141_DO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000ffae5504)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_DO6),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_CO6),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0c0c00000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_B5Q),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y141_SLICE_X5Y141_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05555cccc5555)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_ALUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_AO5),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_DO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033333333)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033a0b30000a0a0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0cfc0cfc0c0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_DO5),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_CO6),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0aaf0aa)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_ALUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaac00c)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_DO6),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaccc8ccc8ccc8)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_DLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_BO6),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0e0e000e000e00)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_BO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaac0aa00)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_DQ),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0aaccccf0aa)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_ALUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_ALUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffdffff)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_DLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I3(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001003300010000)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_CLUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_BO6),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbfffffffeff)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00f3f3c0c0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y138_SLICE_X8Y138_AQ),
.I3(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_DLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001030)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffbff)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefef7f7fffff)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I3(1'b1),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y135_SLICE_X14Y135_AO6),
.Q(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500000045444444)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_DLUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_C5Q),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I5(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffaaff02)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_CLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I2(CLBLM_R_X11Y135_SLICE_X15Y135_DO6),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_DO6),
.I5(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22002200fdfdffff)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb800b8ffb800b8)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_ALUT (
.I0(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100010000000300)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_DLUT (
.I0(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I1(CLBLM_R_X11Y138_SLICE_X15Y138_AO6),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_DO6),
.I3(CLBLM_R_X11Y135_SLICE_X15Y135_CO6),
.I4(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_BO6),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddffddffd0f0ddff)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_CLUT (
.I0(CLBLM_L_X12Y138_SLICE_X16Y138_AO6),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_BO5),
.I3(RIOB33_X105Y143_IOB_X1Y144_I),
.I4(LIOB33_X0Y51_IOB_X0Y52_I),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000abaaefaa)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_BLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_BO6),
.I2(CLBLM_L_X10Y134_SLICE_X13Y134_BQ),
.I3(CLBLM_R_X11Y138_SLICE_X15Y138_BO6),
.I4(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_BO6),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaffaaddd0fff0)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_ALUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.I4(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h004400440f4f0044)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_DLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.I1(LIOB33_X0Y51_IOB_X0Y51_I),
.I2(CLBLM_L_X12Y138_SLICE_X16Y138_BO6),
.I3(CLBLM_R_X11Y135_SLICE_X14Y135_BO5),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00550c5d00000c0c)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_CLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I2(CLBLM_L_X12Y138_SLICE_X16Y138_BO6),
.I3(CLBLM_R_X11Y135_SLICE_X14Y135_BO5),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I5(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000f0000044f4)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X11Y135_SLICE_X14Y135_BO5),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.I5(CLBLM_L_X12Y138_SLICE_X16Y138_BO6),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0f50400040)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_ALUT (
.I0(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I4(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f3f3f1f1)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_DLUT (
.I0(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000300010001)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_CLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_DO6),
.I3(CLBLM_R_X7Y137_SLICE_X9Y137_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y135_SLICE_X15Y135_BO6),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0e1f0e1e1)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_DO6),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_CO6),
.I3(CLBLM_R_X11Y135_SLICE_X15Y135_BO6),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I5(CLBLM_R_X7Y137_SLICE_X9Y137_CO6),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfabbaaf3f03300)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_ALUT (
.I0(CLBLM_R_X11Y138_SLICE_X15Y138_DO6),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I2(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I4(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.Q(CLBLM_R_X11Y137_SLICE_X14Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y137_SLICE_X14Y137_AO6),
.Q(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaaa5556a9a956)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I1(CLBLM_R_X11Y137_SLICE_X15Y137_CO6),
.I2(CLBLM_R_X11Y137_SLICE_X15Y137_DO6),
.I3(CLBLM_L_X10Y138_SLICE_X13Y138_CO6),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_BO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff84ff48ff48ff84)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_CLUT (
.I0(CLBLM_R_X11Y136_SLICE_X15Y136_BO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_AO5),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_DO6),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_DO6),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000005f004f)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_BLUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_CO6),
.I1(CLBLM_L_X12Y138_SLICE_X16Y138_CO6),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_CO6),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X13Y138_CO6),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_CO6),
.I2(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y140_SLICE_X11Y140_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbfffffffa)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_DLUT (
.I0(CLBLM_L_X10Y137_SLICE_X13Y137_AO5),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_DO6),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.I4(CLBLM_R_X7Y137_SLICE_X8Y137_DO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_C5Q),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcfcd0000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_CLUT (
.I0(CLBLM_R_X11Y138_SLICE_X15Y138_CO6),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_CO6),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I3(CLBLM_L_X12Y137_SLICE_X16Y137_DO6),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2322233322222222)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_BLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_CO6),
.I2(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_BO6),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I5(CLBLM_R_X11Y138_SLICE_X15Y138_CO6),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdc)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_ALUT (
.I0(CLBLM_R_X11Y137_SLICE_X15Y137_BO6),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_AO6),
.I5(CLBLM_L_X10Y137_SLICE_X13Y137_BO6),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfefcfefcceeccee)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_DLUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_BO5),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.I3(CLBLM_R_X11Y138_SLICE_X14Y138_AO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_DQ),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_DO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000c555d000c)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_CLUT (
.I0(CLBLM_L_X12Y138_SLICE_X16Y138_BO6),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_DO6),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I4(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_CO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88aa080accff0c0f)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_BLUT (
.I0(CLBLM_R_X11Y139_SLICE_X15Y139_BO6),
.I1(CLBLM_L_X12Y137_SLICE_X16Y137_BO6),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I4(CLBLM_R_X11Y138_SLICE_X14Y138_AO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_BO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbfffffdffff)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_AO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7350735073507350)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_DLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_AO5),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_C5Q),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_DO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033031101)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_CLUT (
.I0(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.I1(CLBLM_R_X11Y138_SLICE_X14Y138_CO6),
.I2(RIOB33_X105Y145_IOB_X1Y145_I),
.I3(CLBLM_R_X11Y138_SLICE_X15Y138_AO5),
.I4(CLBLM_R_X11Y138_SLICE_X14Y138_AO5),
.I5(CLBLM_L_X12Y138_SLICE_X16Y138_AO5),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_CO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00008a8a0000008a)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_BLUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_CO6),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_BO6),
.I5(CLBLM_R_X11Y138_SLICE_X15Y138_AO5),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_BO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c0a0fffffff0)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_AO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X14Y139_AO6),
.Q(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X14Y139_BO6),
.Q(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f300e00020)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_DLUT (
.I0(RIOB33_X105Y141_IOB_X1Y141_I),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_DO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000f0f5f5f5f5f)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_CQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y137_SLICE_X14Y137_BO6),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_CO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfe0efe0e)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_BLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_DQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BO5),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_BO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50fe54fe54)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_AO5),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BO5),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_AO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000020)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I2(CLBLM_R_X3Y139_SLICE_X3Y139_B5Q),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_DO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffbfffaffff)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_CLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_DO6),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_CO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff55ff00004450)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I1(RIOB33_X105Y139_IOB_X1Y139_I),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_BO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffffffffd)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_ALUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_AO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaff00aaaa0000)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y139_IOB_X1Y140_I),
.I4(RIOB33_X105Y141_IOB_X1Y141_I),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_DO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff11ff5fffbbff5f)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_CLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I1(RIOB33_X105Y139_IOB_X1Y140_I),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I4(CLBLL_L_X4Y139_SLICE_X5Y139_D5Q),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_CO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heca0eca03333ffff)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y145_I),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_C5Q),
.I2(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_BO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00a0f5a0f5)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_AO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_AO6),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_DO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefaeeaafcf0cc00)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_CLUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I4(RIOB33_X105Y143_IOB_X1Y144_I),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_CO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefefe)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_BLUT (
.I0(CLBLM_L_X12Y138_SLICE_X16Y138_DO6),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I2(CLBLM_L_X12Y137_SLICE_X17Y137_AO6),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLM_R_X11Y140_SLICE_X15Y140_CO6),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_BO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffeeffcc)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_DO6),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_BQ),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_BO6),
.I4(RIOB33_X105Y139_IOB_X1Y139_I),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_AO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X14Y141_AO6),
.Q(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000800000000)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_DLUT (
.I0(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_BO5),
.I5(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_DO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333133333333333)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_CLUT (
.I0(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_AO6),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_DO5),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_BO5),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_CO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4555ffff0fff0fff)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I2(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_DO6),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_BO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc0caaaaf000)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_ALUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_DQ),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_BO5),
.I2(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I3(CLBLM_R_X11Y141_SLICE_X14Y141_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_DO6),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_AO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X15Y141_AO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X15Y141_BO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_DLUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_DO6),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I3(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I5(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_DO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7ffffffffff)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_CLUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_DO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I3(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I5(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_CO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4a0f5a0a0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_BO6),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.I3(CLBLM_R_X11Y141_SLICE_X14Y141_BO5),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_BO5),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_BO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff001010ff001f1f)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_ALUT (
.I0(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_AO6),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_CO6),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_AO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X18Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X18Y139_DO5),
.O6(CLBLM_R_X13Y139_SLICE_X18Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55f5f5f5f5)
  ) CLBLM_R_X13Y139_SLICE_X18Y139_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_CQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X18Y139_CO5),
.O6(CLBLM_R_X13Y139_SLICE_X18Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffff00ffff)
  ) CLBLM_R_X13Y139_SLICE_X18Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y137_SLICE_X15Y137_AO6),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_CO6),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X18Y139_BO5),
.O6(CLBLM_R_X13Y139_SLICE_X18Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff330f0fffff)
  ) CLBLM_R_X13Y139_SLICE_X18Y139_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I2(CLBLM_R_X11Y136_SLICE_X15Y136_CO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X18Y139_AO5),
.O6(CLBLM_R_X13Y139_SLICE_X18Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_DO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_CO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_BO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y125_IOB_X1Y125_I),
.I2(1'b1),
.I3(RIOB33_X105Y125_IOB_X1Y126_I),
.I4(1'b1),
.I5(RIOB33_X105Y127_IOB_X1Y127_I),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y63_IOB_X0Y64_OBUF (
.I(CLBLM_R_X5Y130_SLICE_X7Y130_AO6),
.O(LIOB33_X0Y63_IOB_X0Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y65_OBUF (
.I(CLBLM_R_X5Y130_SLICE_X7Y130_BO6),
.O(LIOB33_X0Y65_IOB_X0Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y66_OBUF (
.I(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.O(LIOB33_X0Y65_IOB_X0Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLM_R_X5Y130_SLICE_X6Y130_CQ),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLM_R_X3Y139_SLICE_X3Y139_CQ),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X4Y131_SLICE_X5Y131_D5Q),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_A5Q),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(CLBLM_R_X3Y134_SLICE_X3Y134_CQ),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLL_L_X4Y134_SLICE_X4Y134_B5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X6Y138_C5Q),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_R_X7Y129_SLICE_X9Y129_A5Q),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_L_X10Y131_SLICE_X12Y131_C5Q),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X1Y135_CQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X10Y135_SLICE_X12Y135_C5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X1Y135_CQ),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X4Y131_SLICE_X5Y131_DQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X1Y135_CQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X2Y75_SLICE_X0Y75_AO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X2Y137_SLICE_X0Y137_AO5),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X4Y137_SLICE_X4Y137_D5Q),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y138_SLICE_X3Y138_B5Q),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X0Y139_BQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y138_SLICE_X5Y138_CQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X1Y135_CQ),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLM_R_X3Y139_SLICE_X2Y139_DO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLM_R_X5Y142_SLICE_X6Y142_DO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLM_R_X3Y139_SLICE_X2Y139_DO5),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X1Y135_CQ),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(CLBLM_R_X5Y141_SLICE_X6Y141_C5Q),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X1Y135_CQ),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X5Y140_DQ),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X4Y142_CO6),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X5Y140_DO5),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_I),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X0Y139_AQ),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(CLBLM_R_X3Y133_SLICE_X3Y133_DO6),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(CLBLM_R_X3Y165_SLICE_X2Y165_AO6),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(CLBLM_R_X3Y140_SLICE_X2Y140_CO5),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(CLBLL_L_X4Y143_SLICE_X5Y143_DO6),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(1'b1),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLM_R_X3Y140_SLICE_X3Y140_C5Q),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(CLBLM_R_X3Y133_SLICE_X2Y133_DO5),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(1'b1),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_R_X7Y143_SLICE_X8Y143_DO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X7Y138_A5Q),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X7Y138_B5Q),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_L_X10Y141_SLICE_X13Y141_A5Q),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(CLBLM_R_X13Y139_SLICE_X18Y139_AO6),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_L_X8Y143_SLICE_X11Y143_CO6),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X5Y140_DQ),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X5Y140_DO5),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X4Y142_CO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X3Y141_SLICE_X3Y141_DO6),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X3Y140_SLICE_X3Y140_A5Q),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X0Y139_AQ),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(1'b0),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLL_L_X4Y143_SLICE_X5Y143_DO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_L_X8Y143_SLICE_X11Y143_AO6),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X13Y139_SLICE_X18Y139_AO5),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_R_X13Y139_SLICE_X18Y139_CO5),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_L_X12Y139_SLICE_X16Y139_AO6),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_R_X13Y139_SLICE_X18Y139_BO6),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X13Y139_SLICE_X18Y139_CO6),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_L_X12Y139_SLICE_X16Y139_AO5),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y139_SLICE_X17Y139_AO6),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X11Y139_SLICE_X14Y139_CO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X13Y139_SLICE_X18Y139_BO5),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(1'b1),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B = CLBLL_L_X2Y75_SLICE_X0Y75_BO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C = CLBLL_L_X2Y75_SLICE_X0Y75_CO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D = CLBLL_L_X2Y75_SLICE_X0Y75_DO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A = CLBLL_L_X2Y75_SLICE_X1Y75_AO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B = CLBLL_L_X2Y75_SLICE_X1Y75_BO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C = CLBLL_L_X2Y75_SLICE_X1Y75_CO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D = CLBLL_L_X2Y75_SLICE_X1Y75_DO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A = CLBLL_L_X2Y135_SLICE_X0Y135_AO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B = CLBLL_L_X2Y135_SLICE_X0Y135_BO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C = CLBLL_L_X2Y135_SLICE_X0Y135_CO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D = CLBLL_L_X2Y135_SLICE_X0Y135_DO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A = CLBLL_L_X2Y135_SLICE_X1Y135_AO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B = CLBLL_L_X2Y135_SLICE_X1Y135_BO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C = CLBLL_L_X2Y135_SLICE_X1Y135_CO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D = CLBLL_L_X2Y135_SLICE_X1Y135_DO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A = CLBLL_L_X2Y137_SLICE_X0Y137_AO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B = CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C = CLBLL_L_X2Y137_SLICE_X0Y137_CO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D = CLBLL_L_X2Y137_SLICE_X0Y137_DO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_AMUX = CLBLL_L_X2Y137_SLICE_X0Y137_AO5;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A = CLBLL_L_X2Y137_SLICE_X1Y137_AO6;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B = CLBLL_L_X2Y137_SLICE_X1Y137_BO6;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C = CLBLL_L_X2Y137_SLICE_X1Y137_CO6;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D = CLBLL_L_X2Y137_SLICE_X1Y137_DO6;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_CMUX = CLBLL_L_X2Y137_SLICE_X1Y137_C5Q;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B = CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C = CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D = CLBLL_L_X2Y138_SLICE_X0Y138_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A = CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B = CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C = CLBLL_L_X2Y138_SLICE_X1Y138_CO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D = CLBLL_L_X2Y138_SLICE_X1Y138_DO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A = CLBLL_L_X2Y139_SLICE_X0Y139_AO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B = CLBLL_L_X2Y139_SLICE_X0Y139_BO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C = CLBLL_L_X2Y139_SLICE_X0Y139_CO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D = CLBLL_L_X2Y139_SLICE_X0Y139_DO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_BMUX = CLBLL_L_X2Y139_SLICE_X0Y139_B5Q;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A = CLBLL_L_X2Y139_SLICE_X1Y139_AO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B = CLBLL_L_X2Y139_SLICE_X1Y139_BO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C = CLBLL_L_X2Y139_SLICE_X1Y139_CO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D = CLBLL_L_X2Y139_SLICE_X1Y139_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A = CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_CMUX = CLBLL_L_X4Y129_SLICE_X4Y129_CO5;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A = CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C = CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_DMUX = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_AMUX = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_BMUX = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_CMUX = CLBLL_L_X4Y131_SLICE_X4Y131_C5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_DMUX = CLBLL_L_X4Y131_SLICE_X4Y131_DO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B = CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C = CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_CMUX = CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_DMUX = CLBLL_L_X4Y131_SLICE_X5Y131_D5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B = CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C = CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A = CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B = CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D = CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_BMUX = CLBLL_L_X4Y133_SLICE_X4Y133_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_CMUX = CLBLL_L_X4Y133_SLICE_X4Y133_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_DMUX = CLBLL_L_X4Y133_SLICE_X4Y133_D5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A = CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_CMUX = CLBLL_L_X4Y133_SLICE_X5Y133_C5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B = CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_AMUX = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_BMUX = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_CMUX = CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_BMUX = CLBLL_L_X4Y134_SLICE_X5Y134_BO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_DMUX = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A = CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B = CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C = CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D = CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_AMUX = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_BMUX = CLBLL_L_X4Y135_SLICE_X4Y135_B5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_DMUX = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A = CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B = CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C = CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D = CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_AMUX = CLBLL_L_X4Y135_SLICE_X5Y135_A5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_BMUX = CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A = CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B = CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C = CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D = CLBLL_L_X4Y136_SLICE_X4Y136_DO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_AMUX = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_BMUX = CLBLL_L_X4Y136_SLICE_X4Y136_B5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_CMUX = CLBLL_L_X4Y136_SLICE_X4Y136_C5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_DMUX = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A = CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D = CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_BMUX = CLBLL_L_X4Y136_SLICE_X5Y136_B5Q;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_CMUX = CLBLL_L_X4Y136_SLICE_X5Y136_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B = CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C = CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D = CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_CMUX = CLBLL_L_X4Y137_SLICE_X4Y137_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_DMUX = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A = CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B = CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C = CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D = CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_CMUX = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_DMUX = CLBLL_L_X4Y137_SLICE_X5Y137_D5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D = CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A = CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B = CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C = CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_AMUX = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_BMUX = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_CMUX = CLBLL_L_X4Y138_SLICE_X5Y138_C5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A = CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C = CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D = CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_AMUX = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_CMUX = CLBLL_L_X4Y139_SLICE_X4Y139_C5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A = CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B = CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C = CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D = CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_CMUX = CLBLL_L_X4Y139_SLICE_X5Y139_C5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_DMUX = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_CMUX = CLBLL_L_X4Y140_SLICE_X4Y140_C5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_AMUX = CLBLL_L_X4Y140_SLICE_X5Y140_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_BMUX = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_CMUX = CLBLL_L_X4Y140_SLICE_X5Y140_C5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_DMUX = CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A = CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B = CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_CMUX = CLBLL_L_X4Y141_SLICE_X4Y141_C5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A = CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_CMUX = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A = CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_AMUX = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_CMUX = CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A = CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D = CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_AMUX = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_BMUX = CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_CMUX = CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_BMUX = CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CMUX = CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A = CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C = CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_DMUX = CLBLM_L_X8Y131_SLICE_X10Y131_D5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A = CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_AMUX = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CMUX = CLBLM_L_X8Y131_SLICE_X11Y131_C5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A = CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_AMUX = CLBLM_L_X8Y132_SLICE_X10Y132_A5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_CMUX = CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_BMUX = CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_CMUX = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_AMUX = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A = CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B = CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_AMUX = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_BMUX = CLBLM_L_X8Y134_SLICE_X10Y134_B5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A = CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B = CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_DMUX = CLBLM_L_X8Y134_SLICE_X11Y134_DO5;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A = CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_AMUX = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A = CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_BMUX = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A = CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_DMUX = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A = CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B = CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A = CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B = CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C = CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D = CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A = CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B = CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D = CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C = CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A = CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_BMUX = CLBLM_L_X8Y138_SLICE_X11Y138_BO5;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A = CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C = CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D = CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_BMUX = CLBLM_L_X8Y139_SLICE_X10Y139_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_CMUX = CLBLM_L_X8Y139_SLICE_X10Y139_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A = CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B = CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_CMUX = CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_DMUX = CLBLM_L_X8Y139_SLICE_X11Y139_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A = CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B = CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_BMUX = CLBLM_L_X8Y140_SLICE_X10Y140_B5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_CMUX = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_DMUX = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_CMUX = CLBLM_L_X8Y140_SLICE_X11Y140_C5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B = CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A = CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C = CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A = CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_AMUX = CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A = CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_CMUX = CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CMUX = CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_CMUX = CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A = CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_AMUX = CLBLM_L_X10Y133_SLICE_X12Y133_A5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A = CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_DMUX = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A = CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B = CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D = CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_BMUX = CLBLM_L_X10Y134_SLICE_X12Y134_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_DMUX = CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A = CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_CMUX = CLBLM_L_X10Y134_SLICE_X13Y134_C5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B = CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_CMUX = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_AMUX = CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_BMUX = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A = CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_AMUX = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CMUX = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_AMUX = CLBLM_L_X10Y137_SLICE_X12Y137_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_BMUX = CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_CMUX = CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A = CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_AMUX = CLBLM_L_X10Y137_SLICE_X13Y137_AO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_CMUX = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_BMUX = CLBLM_L_X10Y138_SLICE_X12Y138_B5Q;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_CMUX = CLBLM_L_X10Y138_SLICE_X12Y138_C5Q;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A = CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B = CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C = CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D = CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A = CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D = CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_AMUX = CLBLM_L_X10Y139_SLICE_X12Y139_AO5;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_BMUX = CLBLM_L_X10Y139_SLICE_X12Y139_BO5;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_CMUX = CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A = CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C = CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D = CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_AMUX = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_BMUX = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_CMUX = CLBLM_L_X10Y139_SLICE_X13Y139_C5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A = CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B = CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_AMUX = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_BMUX = CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_CMUX = CLBLM_L_X10Y140_SLICE_X12Y140_C5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_DMUX = CLBLM_L_X10Y140_SLICE_X12Y140_DO5;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A = CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B = CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C = CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_AMUX = CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_BMUX = CLBLM_L_X10Y140_SLICE_X13Y140_BO5;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_CMUX = CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A = CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C = CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A = CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B = CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_AMUX = CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_CMUX = CLBLM_L_X10Y141_SLICE_X13Y141_CO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_AMUX = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A = CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_DMUX = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_CMUX = CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B = CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C = CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D = CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D = CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C = CLBLM_L_X12Y136_SLICE_X16Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D = CLBLM_L_X12Y136_SLICE_X16Y136_DO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_AMUX = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A = CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C = CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D = CLBLM_L_X12Y136_SLICE_X17Y136_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B = CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_AMUX = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_BMUX = CLBLM_L_X12Y137_SLICE_X16Y137_BO5;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A = CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B = CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C = CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A = CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B = CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C = CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D = CLBLM_L_X12Y138_SLICE_X16Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_AMUX = CLBLM_L_X12Y138_SLICE_X16Y138_AO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_BMUX = CLBLM_L_X12Y138_SLICE_X16Y138_BO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_CMUX = CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A = CLBLM_L_X12Y138_SLICE_X17Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C = CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B = CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C = CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D = CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_AMUX = CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B = CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C = CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B = CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D = CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A = CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B = CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_AMUX = CLBLM_R_X3Y129_SLICE_X3Y129_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_BMUX = CLBLM_R_X3Y129_SLICE_X3Y129_BO5;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B = CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A = CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_DMUX = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A = CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B = CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_AMUX = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A = CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B = CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C = CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D = CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_AMUX = CLBLM_R_X3Y132_SLICE_X3Y132_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_BMUX = CLBLM_R_X3Y132_SLICE_X3Y132_BO5;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A = CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B = CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C = CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D = CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_BMUX = CLBLM_R_X3Y133_SLICE_X2Y133_B5Q;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_CMUX = CLBLM_R_X3Y133_SLICE_X2Y133_C5Q;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_DMUX = CLBLM_R_X3Y133_SLICE_X2Y133_DO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_BMUX = CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A = CLBLM_R_X3Y134_SLICE_X2Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B = CLBLM_R_X3Y134_SLICE_X2Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C = CLBLM_R_X3Y134_SLICE_X2Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D = CLBLM_R_X3Y134_SLICE_X2Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_AMUX = CLBLM_R_X3Y134_SLICE_X2Y134_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A = CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B = CLBLM_R_X3Y134_SLICE_X3Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C = CLBLM_R_X3Y134_SLICE_X3Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_CMUX = CLBLM_R_X3Y134_SLICE_X3Y134_C5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_DMUX = CLBLM_R_X3Y134_SLICE_X3Y134_D5Q;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A = CLBLM_R_X3Y135_SLICE_X2Y135_AO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B = CLBLM_R_X3Y135_SLICE_X2Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C = CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D = CLBLM_R_X3Y135_SLICE_X2Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_AMUX = CLBLM_R_X3Y135_SLICE_X2Y135_AO5;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_BMUX = CLBLM_R_X3Y135_SLICE_X2Y135_BO5;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A = CLBLM_R_X3Y135_SLICE_X3Y135_AO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B = CLBLM_R_X3Y135_SLICE_X3Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C = CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D = CLBLM_R_X3Y135_SLICE_X3Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_CMUX = CLBLM_R_X3Y135_SLICE_X3Y135_C5Q;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A = CLBLM_R_X3Y136_SLICE_X2Y136_AO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B = CLBLM_R_X3Y136_SLICE_X2Y136_BO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C = CLBLM_R_X3Y136_SLICE_X2Y136_CO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D = CLBLM_R_X3Y136_SLICE_X2Y136_DO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_DMUX = CLBLM_R_X3Y136_SLICE_X2Y136_DO5;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A = CLBLM_R_X3Y136_SLICE_X3Y136_AO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B = CLBLM_R_X3Y136_SLICE_X3Y136_BO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C = CLBLM_R_X3Y136_SLICE_X3Y136_CO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D = CLBLM_R_X3Y136_SLICE_X3Y136_DO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_AMUX = CLBLM_R_X3Y136_SLICE_X3Y136_A5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_BMUX = CLBLM_R_X3Y136_SLICE_X3Y136_B5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_CMUX = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_DMUX = CLBLM_R_X3Y136_SLICE_X3Y136_D5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A = CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B = CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C = CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D = CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_DMUX = CLBLM_R_X3Y137_SLICE_X2Y137_D5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A = CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B = CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C = CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D = CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_BMUX = CLBLM_R_X3Y137_SLICE_X3Y137_B5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_CMUX = CLBLM_R_X3Y137_SLICE_X3Y137_C5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_DMUX = CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A = CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B = CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C = CLBLM_R_X3Y138_SLICE_X2Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D = CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_AMUX = CLBLM_R_X3Y138_SLICE_X2Y138_A5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A = CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B = CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C = CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D = CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_AMUX = CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_BMUX = CLBLM_R_X3Y138_SLICE_X3Y138_B5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_CMUX = CLBLM_R_X3Y138_SLICE_X3Y138_C5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_DMUX = CLBLM_R_X3Y138_SLICE_X3Y138_D5Q;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A = CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B = CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C = CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D = CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_AMUX = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_BMUX = CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_CMUX = CLBLM_R_X3Y139_SLICE_X2Y139_CO5;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_DMUX = CLBLM_R_X3Y139_SLICE_X2Y139_DO5;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A = CLBLM_R_X3Y139_SLICE_X3Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C = CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D = CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_AMUX = CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_BMUX = CLBLM_R_X3Y139_SLICE_X3Y139_B5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_CMUX = CLBLM_R_X3Y139_SLICE_X3Y139_C5Q;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A = CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B = CLBLM_R_X3Y140_SLICE_X2Y140_BO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C = CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_AMUX = CLBLM_R_X3Y140_SLICE_X2Y140_A5Q;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_CMUX = CLBLM_R_X3Y140_SLICE_X2Y140_CO5;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A = CLBLM_R_X3Y140_SLICE_X3Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B = CLBLM_R_X3Y140_SLICE_X3Y140_BO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C = CLBLM_R_X3Y140_SLICE_X3Y140_CO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D = CLBLM_R_X3Y140_SLICE_X3Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_AMUX = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_CMUX = CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_DMUX = CLBLM_R_X3Y140_SLICE_X3Y140_DO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D = CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C = CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_A = CLBLM_R_X3Y165_SLICE_X2Y165_AO6;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_B = CLBLM_R_X3Y165_SLICE_X2Y165_BO6;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_C = CLBLM_R_X3Y165_SLICE_X2Y165_CO6;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_D = CLBLM_R_X3Y165_SLICE_X2Y165_DO6;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_A = CLBLM_R_X3Y165_SLICE_X3Y165_AO6;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_B = CLBLM_R_X3Y165_SLICE_X3Y165_BO6;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_C = CLBLM_R_X3Y165_SLICE_X3Y165_CO6;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_D = CLBLM_R_X3Y165_SLICE_X3Y165_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CMUX = CLBLM_R_X5Y130_SLICE_X6Y130_C5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A = CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B = CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CMUX = CLBLM_R_X5Y131_SLICE_X6Y131_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_DMUX = CLBLM_R_X5Y131_SLICE_X6Y131_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A = CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B = CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C = CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B = CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_AMUX = CLBLM_R_X5Y132_SLICE_X6Y132_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_DMUX = CLBLM_R_X5Y132_SLICE_X6Y132_DO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A = CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A = CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A = CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_AMUX = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_BMUX = CLBLM_R_X5Y133_SLICE_X7Y133_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_CMUX = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_DMUX = CLBLM_R_X5Y133_SLICE_X7Y133_D5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_BMUX = CLBLM_R_X5Y134_SLICE_X6Y134_B5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_CMUX = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A = CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C = CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_CMUX = CLBLM_R_X5Y134_SLICE_X7Y134_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_DMUX = CLBLM_R_X5Y134_SLICE_X7Y134_D5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A = CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B = CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_CMUX = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_DMUX = CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A = CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_BMUX = CLBLM_R_X5Y135_SLICE_X7Y135_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A = CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B = CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_BMUX = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_CMUX = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_DMUX = CLBLM_R_X5Y136_SLICE_X6Y136_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B = CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C = CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_AMUX = CLBLM_R_X5Y136_SLICE_X7Y136_A5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_BMUX = CLBLM_R_X5Y136_SLICE_X7Y136_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_CMUX = CLBLM_R_X5Y136_SLICE_X7Y136_C5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B = CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_BMUX = CLBLM_R_X5Y137_SLICE_X6Y137_B5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_CMUX = CLBLM_R_X5Y137_SLICE_X6Y137_C5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_DMUX = CLBLM_R_X5Y137_SLICE_X6Y137_D5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A = CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B = CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C = CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_CMUX = CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C = CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_BMUX = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_CMUX = CLBLM_R_X5Y138_SLICE_X6Y138_C5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A = CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B = CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_AMUX = CLBLM_R_X5Y138_SLICE_X7Y138_A5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_BMUX = CLBLM_R_X5Y138_SLICE_X7Y138_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_CMUX = CLBLM_R_X5Y138_SLICE_X7Y138_C5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A = CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C = CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_AMUX = CLBLM_R_X5Y139_SLICE_X6Y139_A5Q;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A = CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B = CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C = CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_AMUX = CLBLM_R_X5Y139_SLICE_X7Y139_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_AMUX = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_BMUX = CLBLM_R_X5Y140_SLICE_X6Y140_B5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_CMUX = CLBLM_R_X5Y140_SLICE_X6Y140_C5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A = CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B = CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C = CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_BMUX = CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_CMUX = CLBLM_R_X5Y140_SLICE_X7Y140_C5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_DMUX = CLBLM_R_X5Y140_SLICE_X7Y140_D5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A = CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B = CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C = CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_BMUX = CLBLM_R_X5Y141_SLICE_X6Y141_B5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_CMUX = CLBLM_R_X5Y141_SLICE_X6Y141_C5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_DMUX = CLBLM_R_X5Y141_SLICE_X6Y141_DO5;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B = CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C = CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_CMUX = CLBLM_R_X5Y141_SLICE_X7Y141_CO5;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A = CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B = CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A = CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_CMUX = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_DMUX = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C = CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D = CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_AMUX = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A = CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_CMUX = CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_DMUX = CLBLM_R_X5Y143_SLICE_X7Y143_DO5;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A = CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C = CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A = CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C = CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_AMUX = CLBLM_R_X5Y144_SLICE_X7Y144_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A = CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B = CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A = CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_AMUX = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A = CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B = CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CMUX = CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_DMUX = CLBLM_R_X7Y130_SLICE_X8Y130_DO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A = CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_BMUX = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CMUX = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CMUX = CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A = CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_AMUX = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_BMUX = CLBLM_R_X7Y131_SLICE_X9Y131_B5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CMUX = CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A = CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_BMUX = CLBLM_R_X7Y132_SLICE_X8Y132_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_CMUX = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_AMUX = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A = CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B = CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C = CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_AMUX = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_DMUX = CLBLM_R_X7Y133_SLICE_X8Y133_DO5;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A = CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C = CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_AMUX = CLBLM_R_X7Y133_SLICE_X9Y133_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_BMUX = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_CMUX = CLBLM_R_X7Y133_SLICE_X9Y133_CO5;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A = CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B = CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C = CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_DMUX = CLBLM_R_X7Y134_SLICE_X8Y134_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A = CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B = CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C = CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_BMUX = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_DMUX = CLBLM_R_X7Y134_SLICE_X9Y134_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A = CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A = CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B = CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_AMUX = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_BMUX = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A = CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B = CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_AMUX = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_BMUX = CLBLM_R_X7Y136_SLICE_X8Y136_B5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_DMUX = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A = CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_CMUX = CLBLM_R_X7Y136_SLICE_X9Y136_C5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B = CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C = CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_BMUX = CLBLM_R_X7Y137_SLICE_X8Y137_B5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_CMUX = CLBLM_R_X7Y137_SLICE_X8Y137_C5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A = CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B = CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_AMUX = CLBLM_R_X7Y137_SLICE_X9Y137_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A = CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B = CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C = CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D = CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_AMUX = CLBLM_R_X7Y138_SLICE_X8Y138_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A = CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C = CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B = CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A = CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_AMUX = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A = CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B = CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C = CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_BMUX = CLBLM_R_X7Y140_SLICE_X8Y140_B5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_DMUX = CLBLM_R_X7Y140_SLICE_X8Y140_D5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A = CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B = CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C = CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_CMUX = CLBLM_R_X7Y140_SLICE_X9Y140_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_DMUX = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A = CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_AMUX = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_DMUX = CLBLM_R_X7Y141_SLICE_X8Y141_DO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C = CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D = CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_CMUX = CLBLM_R_X7Y141_SLICE_X9Y141_C5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_DMUX = CLBLM_R_X7Y141_SLICE_X9Y141_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A = CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_AMUX = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_CMUX = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B = CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_CMUX = CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A = CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C = CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_AMUX = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_BMUX = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_DMUX = CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A = CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B = CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C = CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_AMUX = CLBLM_R_X7Y143_SLICE_X9Y143_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_BMUX = CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A = CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_DMUX = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B = CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C = CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D = CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_AMUX = CLBLM_R_X11Y134_SLICE_X14Y134_A5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_BMUX = CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_AMUX = CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D = CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_BMUX = CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B = CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C = CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D = CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_AMUX = CLBLM_R_X11Y136_SLICE_X14Y136_AO5;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B = CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_AMUX = CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_AMUX = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_BMUX = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C = CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D = CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_BMUX = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A = CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B = CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C = CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D = CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_AMUX = CLBLM_R_X11Y138_SLICE_X14Y138_AO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A = CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B = CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_AMUX = CLBLM_R_X11Y138_SLICE_X15Y138_AO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A = CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B = CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C = CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_CMUX = CLBLM_R_X11Y139_SLICE_X14Y139_CO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_DMUX = CLBLM_R_X11Y139_SLICE_X14Y139_DO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B = CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_AMUX = CLBLM_R_X11Y139_SLICE_X15Y139_AO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_BMUX = CLBLM_R_X11Y139_SLICE_X15Y139_BO5;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D = CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_AMUX = CLBLM_R_X11Y140_SLICE_X14Y140_AO5;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_BMUX = CLBLM_R_X11Y140_SLICE_X14Y140_BO5;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_DMUX = CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A = CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B = CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C = CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D = CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A = CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B = CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_BMUX = CLBLM_R_X11Y141_SLICE_X14Y141_BO5;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A = CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B = CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C = CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A = CLBLM_R_X13Y139_SLICE_X18Y139_AO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C = CLBLM_R_X13Y139_SLICE_X18Y139_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D = CLBLM_R_X13Y139_SLICE_X18Y139_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_AMUX = CLBLM_R_X13Y139_SLICE_X18Y139_AO5;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_BMUX = CLBLM_R_X13Y139_SLICE_X18Y139_BO5;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_CMUX = CLBLM_R_X13Y139_SLICE_X18Y139_CO5;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C = CLBLM_R_X13Y139_SLICE_X19Y139_CO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A = CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B = CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C = CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D = CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B = CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C = CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D = CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_OQ = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_TQ = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_OQ = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_TQ = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLM_R_X3Y139_SLICE_X3Y139_CQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X5Y138_SLICE_X6Y138_C5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X2Y137_SLICE_X0Y137_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y138_SLICE_X5Y138_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X2Y139_SLICE_X0Y139_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLM_R_X3Y139_SLICE_X2Y139_DO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = CLBLM_R_X5Y141_SLICE_X6Y141_C5Q;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = CLBLL_L_X2Y139_SLICE_X0Y139_AQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = CLBLM_R_X3Y140_SLICE_X2Y140_CO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = CLBLM_R_X3Y133_SLICE_X2Y133_DO5;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_A5Q;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X4Y131_SLICE_X5Y131_D5Q;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = CLBLM_R_X3Y165_SLICE_X2Y165_AO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y138_SLICE_X3Y138_B5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_R_X5Y138_SLICE_X7Y138_A5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = CLBLM_R_X13Y139_SLICE_X18Y139_AO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLL_L_X2Y139_SLICE_X0Y139_AQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = 1'b0;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X13Y139_SLICE_X18Y139_AO5;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_R_X13Y139_SLICE_X18Y139_CO5;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X13Y139_SLICE_X18Y139_BO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X11Y139_SLICE_X14Y139_CO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X13Y139_SLICE_X18Y139_CO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_R_X5Y138_SLICE_X7Y138_B5Q;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLM_R_X3Y139_SLICE_X2Y139_DO5;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C2 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A2 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A4 = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A5 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A6 = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C4 = CLBLM_L_X8Y140_SLICE_X11Y140_DQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_AX = CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C5 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B1 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B3 = CLBLM_R_X7Y134_SLICE_X8Y134_DQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B6 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C6 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C1 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C2 = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C3 = CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C5 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C6 = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D2 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D4 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D6 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A1 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A2 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A4 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A5 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A6 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_AX = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B1 = CLBLM_L_X8Y131_SLICE_X11Y131_C5Q;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B2 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B3 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B4 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B5 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D1 = CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_BX = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D2 = CLBLL_L_X4Y136_SLICE_X5Y136_B5Q;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C1 = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C2 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C3 = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C6 = CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CX = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D1 = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D3 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D6 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A1 = CLBLL_L_X2Y139_SLICE_X0Y139_B5Q;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A2 = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A3 = CLBLL_L_X2Y138_SLICE_X1Y138_AQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A4 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A6 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D4 = CLBLM_R_X11Y138_SLICE_X14Y138_AO5;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B2 = CLBLL_L_X2Y138_SLICE_X1Y138_BQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B3 = CLBLL_L_X2Y138_SLICE_X1Y138_AQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B4 = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B5 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B6 = CLBLM_R_X3Y138_SLICE_X3Y138_B5Q;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D6 = CLBLM_L_X10Y138_SLICE_X12Y138_DQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C3 = CLBLL_L_X4Y139_SLICE_X5Y139_C5Q;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = 1'b1;
  assign LIOB33_X0Y151_IOB_X0Y152_O = CLBLM_R_X5Y141_SLICE_X6Y141_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B6 = 1'b1;
  assign LIOB33_X0Y151_IOB_X0Y151_O = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D4 = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C6 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A3 = CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B1 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D2 = CLBLM_R_X7Y132_SLICE_X8Y132_B5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B2 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B3 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B4 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D3 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A3 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A6 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D4 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D5 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B2 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B6 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D4 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A1 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A2 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A3 = CLBLM_L_X8Y139_SLICE_X11Y139_D5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A5 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A6 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B1 = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B2 = CLBLM_R_X5Y139_SLICE_X7Y139_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B4 = CLBLM_R_X7Y140_SLICE_X8Y140_CQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B5 = CLBLM_R_X7Y136_SLICE_X9Y136_C5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A1 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A3 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A4 = CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A5 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C1 = CLBLM_R_X7Y137_SLICE_X8Y137_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C2 = CLBLM_R_X7Y140_SLICE_X8Y140_CQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B1 = CLBLM_R_X5Y131_SLICE_X6Y131_DQ;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A1 = CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A3 = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A5 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B3 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B4 = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B1 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B2 = CLBLL_L_X4Y139_SLICE_X4Y139_C5Q;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B3 = CLBLL_L_X2Y139_SLICE_X0Y139_AQ;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B5 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C2 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D6 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A1 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A2 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A3 = CLBLM_R_X3Y138_SLICE_X2Y138_DQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A5 = CLBLL_L_X2Y137_SLICE_X0Y137_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A6 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B1 = CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B2 = CLBLL_L_X2Y139_SLICE_X1Y139_BQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B3 = CLBLL_L_X2Y137_SLICE_X1Y137_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B4 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B6 = CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C1 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C2 = CLBLL_L_X2Y139_SLICE_X1Y139_CQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C4 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C5 = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C6 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y153_IOB_X0Y153_O = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign LIOB33_X0Y153_IOB_X0Y154_O = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D2 = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D3 = CLBLL_L_X2Y139_SLICE_X1Y139_DQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D4 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D6 = CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D2 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A1 = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A2 = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A3 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A4 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A5 = CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B1 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B2 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B5 = CLBLL_L_X4Y136_SLICE_X5Y136_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B6 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A1 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A2 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A3 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C1 = CLBLM_L_X10Y140_SLICE_X12Y140_C5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C3 = CLBLM_R_X7Y140_SLICE_X8Y140_DQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B1 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B2 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B3 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B4 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C1 = CLBLM_R_X5Y134_SLICE_X7Y134_DQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C2 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C3 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C5 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D3 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A1 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A2 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A5 = CLBLM_R_X5Y141_SLICE_X7Y141_CO5;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A6 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D2 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D4 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_AX = CLBLM_R_X7Y141_SLICE_X8Y141_DO5;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B1 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B2 = CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B3 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B4 = CLBLM_R_X5Y139_SLICE_X7Y139_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B5 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A2 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A3 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A5 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C2 = CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C3 = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B1 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B2 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B3 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B4 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D1 = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C1 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C2 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C5 = CLBLM_R_X5Y131_SLICE_X6Y131_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D3 = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D4 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D5 = CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D1 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D3 = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D4 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D5 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign LIOB33_X0Y155_IOB_X0Y155_O = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C3 = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X13Y139_SLICE_X18Y139_CO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C2 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C3 = CLBLM_R_X3Y134_SLICE_X3Y134_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A1 = CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A2 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A3 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A4 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A6 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D2 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B1 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B2 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B4 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B6 = CLBLL_L_X4Y136_SLICE_X5Y136_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A2 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A3 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A6 = CLBLL_L_X4Y136_SLICE_X4Y136_B5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C2 = CLBLM_L_X8Y140_SLICE_X11Y140_DQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C3 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B2 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B3 = CLBLM_R_X5Y136_SLICE_X7Y136_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B4 = CLBLL_L_X4Y133_SLICE_X4Y133_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B5 = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B6 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D1 = CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C1 = CLBLM_R_X3Y133_SLICE_X2Y133_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C2 = CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C3 = CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C4 = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C5 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D3 = CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D4 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A1 = CLBLM_R_X7Y139_SLICE_X8Y139_CQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A2 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A4 = CLBLM_R_X3Y140_SLICE_X2Y140_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D1 = CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D2 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D3 = CLBLM_R_X5Y140_SLICE_X7Y140_DQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D4 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D6 = CLBLL_L_X4Y131_SLICE_X5Y131_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B1 = CLBLM_R_X7Y133_SLICE_X9Y133_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A2 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A3 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A4 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A6 = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_AX = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B1 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B2 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B4 = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B5 = CLBLM_R_X5Y134_SLICE_X6Y134_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B1 = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C2 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C3 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C5 = CLBLM_R_X5Y132_SLICE_X6Y132_DO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C6 = CLBLM_R_X3Y135_SLICE_X2Y135_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D2 = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D6 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D1 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D3 = CLBLM_R_X7Y131_SLICE_X9Y131_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D4 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D5 = CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D6 = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D2 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D3 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A6 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A1 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A2 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A3 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A5 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B2 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B4 = CLBLM_R_X5Y143_SLICE_X7Y143_DO5;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B5 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B6 = CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_BX = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A2 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A3 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A5 = CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C2 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C3 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B1 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B2 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B4 = CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B5 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C1 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C3 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C4 = CLBLM_R_X3Y133_SLICE_X2Y133_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C5 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A1 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A2 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A3 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D1 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D3 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D4 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B5 = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B1 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A1 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A3 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A4 = CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A5 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C1 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C2 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B1 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B2 = CLBLM_R_X5Y134_SLICE_X7Y134_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B4 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B5 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B6 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C2 = CLBLM_R_X5Y133_SLICE_X6Y133_CQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C3 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C4 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C5 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C6 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D2 = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D1 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D2 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D3 = CLBLM_R_X5Y133_SLICE_X6Y133_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D4 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C5 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D4 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1 = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A1 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A4 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B1 = CLBLL_L_X4Y139_SLICE_X5Y139_DQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B3 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C4 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B6 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C5 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A1 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A2 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A3 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A6 = CLBLM_R_X5Y136_SLICE_X7Y136_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C1 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C2 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B1 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B2 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B3 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B4 = CLBLM_R_X5Y134_SLICE_X7Y134_D5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B5 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D1 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C2 = CLBLM_R_X3Y133_SLICE_X2Y133_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C3 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C5 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D3 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D4 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A3 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D2 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D3 = CLBLM_R_X5Y136_SLICE_X7Y136_B5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D4 = CLBLM_R_X3Y138_SLICE_X2Y138_DQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D5 = CLBLM_R_X7Y140_SLICE_X9Y140_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A2 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A3 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A4 = CLBLM_R_X5Y133_SLICE_X7Y133_D5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A6 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B1 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B3 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B4 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B5 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D2 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C1 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C4 = CLBLL_L_X2Y135_SLICE_X1Y135_DQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C5 = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D2 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D3 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D4 = CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D5 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D6 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D1 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D2 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D3 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D4 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D5 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C4 = CLBLM_R_X5Y139_SLICE_X6Y139_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B2 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C4 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C6 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C2 = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C3 = CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C6 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A1 = CLBLM_R_X5Y133_SLICE_X6Y133_DQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A2 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A3 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A4 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A6 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign LIOB33_X0Y163_IOB_X0Y163_O = CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B1 = CLBLM_R_X7Y143_SLICE_X9Y143_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B2 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B4 = CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B5 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C1 = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C2 = CLBLL_L_X2Y135_SLICE_X1Y135_DQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C3 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C4 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C5 = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C6 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D1 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D2 = CLBLM_R_X7Y143_SLICE_X9Y143_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D3 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D4 = CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D5 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A2 = CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A3 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A5 = CLBLL_L_X2Y135_SLICE_X1Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A6 = CLBLM_R_X7Y133_SLICE_X9Y133_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B1 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B2 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B4 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B5 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B6 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C2 = CLBLL_L_X4Y135_SLICE_X5Y135_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C3 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C4 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C5 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D1 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D3 = CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D4 = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D5 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D6 = 1'b1;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A1 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A2 = CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A4 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A5 = CLBLM_R_X5Y140_SLICE_X6Y140_C5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B1 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B2 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B4 = CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B5 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C2 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C3 = CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D1 = CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D2 = CLBLM_R_X5Y133_SLICE_X6Y133_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D4 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D5 = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D6 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLM_R_X3Y139_SLICE_X3Y139_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A3 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A4 = CLBLL_L_X4Y137_SLICE_X5Y137_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B1 = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B2 = CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B3 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B4 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C1 = CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C2 = CLBLM_R_X5Y136_SLICE_X6Y136_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C3 = CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C4 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D2 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D4 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A1 = CLBLM_R_X7Y140_SLICE_X9Y140_DQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A2 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A3 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A4 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A6 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B1 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B2 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B4 = CLBLL_L_X2Y137_SLICE_X1Y137_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B5 = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B6 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C1 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C3 = CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C4 = CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D1 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D2 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D3 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D5 = CLBLM_R_X7Y132_SLICE_X8Y132_B5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A2 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A3 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A4 = CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A5 = CLBLM_R_X5Y131_SLICE_X6Y131_DQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A6 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B2 = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B3 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B4 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B5 = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C1 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C2 = CLBLM_R_X5Y133_SLICE_X6Y133_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C3 = CLBLL_L_X4Y135_SLICE_X4Y135_B5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C4 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D2 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D3 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D4 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D5 = CLBLL_L_X4Y133_SLICE_X4Y133_C5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A1 = CLBLM_R_X5Y138_SLICE_X7Y138_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A2 = CLBLM_R_X5Y135_SLICE_X6Y135_DQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A4 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A5 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B1 = CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B3 = CLBLM_R_X5Y136_SLICE_X7Y136_C5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B4 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B5 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B6 = 1'b1;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C2 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C3 = CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C4 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C5 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D1 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D2 = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D3 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D5 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A1 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A2 = CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A3 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A5 = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A6 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B1 = CLBLM_R_X7Y134_SLICE_X9Y134_D5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B2 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B3 = CLBLL_L_X4Y138_SLICE_X5Y138_CQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B5 = CLBLM_R_X5Y138_SLICE_X6Y138_C5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C1 = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C3 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C4 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C5 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D1 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D2 = CLBLM_R_X5Y134_SLICE_X6Y134_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D3 = CLBLM_R_X5Y138_SLICE_X7Y138_CQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D4 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C4 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C5 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C6 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign LIOB33_X0Y171_IOB_X0Y172_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y171_IOB_X0Y171_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D2 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D5 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A1 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A2 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A4 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A5 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C4 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C5 = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B1 = CLBLM_R_X11Y140_SLICE_X14Y140_BO5;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B2 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B3 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B4 = CLBLL_L_X4Y141_SLICE_X4Y141_C5Q;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A3 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A4 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A6 = CLBLM_R_X3Y138_SLICE_X2Y138_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C2 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_AX = CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C3 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B1 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B2 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B3 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B5 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D1 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D3 = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D4 = CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A1 = CLBLM_R_X5Y137_SLICE_X6Y137_DQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A2 = CLBLM_R_X7Y138_SLICE_X8Y138_A5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A3 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A4 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B1 = CLBLM_R_X5Y132_SLICE_X6Y132_A5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B3 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B4 = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A3 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C3 = CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C4 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C5 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D1 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D2 = CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D3 = CLBLM_L_X8Y139_SLICE_X10Y139_B5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D4 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D5 = CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D6 = CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C5 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A1 = CLBLM_R_X7Y141_SLICE_X9Y141_D5Q;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D1 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B1 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B2 = CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D4 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B3 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign LIOB33_X0Y173_IOB_X0Y173_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOB33_X0Y173_IOB_X0Y174_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D5 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D6 = CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B5 = CLBLM_R_X7Y141_SLICE_X9Y141_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C5 = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C6 = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C3 = CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C5 = CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A3 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A4 = CLBLM_R_X5Y137_SLICE_X6Y137_DQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A5 = CLBLM_R_X5Y140_SLICE_X7Y140_C5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B1 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B2 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B3 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C1 = CLBLL_L_X4Y141_SLICE_X4Y141_C5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C2 = CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C3 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C4 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D5 = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D2 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D3 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D4 = CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D5 = CLBLM_R_X5Y138_SLICE_X6Y138_C5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A2 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A3 = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A4 = CLBLM_R_X7Y140_SLICE_X8Y140_D5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B1 = CLBLL_L_X4Y137_SLICE_X4Y137_DQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B4 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B5 = CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B6 = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C2 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C3 = CLBLL_L_X4Y140_SLICE_X4Y140_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C4 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D2 = CLBLM_L_X8Y134_SLICE_X10Y134_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D3 = CLBLL_L_X4Y140_SLICE_X5Y140_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D4 = CLBLM_R_X7Y140_SLICE_X8Y140_D5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D5 = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D6 = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D5 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D2 = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y138_SLICE_X3Y138_B5Q;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A1 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A2 = CLBLM_R_X5Y138_SLICE_X7Y138_CQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A3 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A5 = CLBLM_R_X5Y141_SLICE_X7Y141_CO5;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B1 = CLBLM_R_X5Y140_SLICE_X7Y140_DQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B2 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B3 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B6 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A1 = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A2 = CLBLM_R_X5Y131_SLICE_X6Y131_D5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C4 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C5 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A4 = CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A5 = CLBLL_L_X4Y133_SLICE_X5Y133_C5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A6 = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C1 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B1 = CLBLM_R_X3Y132_SLICE_X3Y132_BO5;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B2 = CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B4 = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B5 = CLBLM_R_X5Y131_SLICE_X6Y131_D5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B6 = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D1 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C1 = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C2 = CLBLL_L_X4Y131_SLICE_X5Y131_D5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C3 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C4 = CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C5 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C6 = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D4 = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A1 = CLBLM_R_X5Y141_SLICE_X6Y141_DO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A3 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A4 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A5 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A6 = CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D2 = CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D4 = CLBLM_R_X3Y132_SLICE_X3Y132_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D5 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D6 = CLBLM_R_X3Y133_SLICE_X2Y133_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B3 = CLBLM_R_X3Y139_SLICE_X3Y139_C5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B4 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B5 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A2 = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A3 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A4 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A5 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A6 = CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C1 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C2 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B4 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B6 = CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D1 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D3 = CLBLM_L_X10Y139_SLICE_X13Y139_C5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D4 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D5 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C6 = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D6 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A4 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A5 = CLBLM_R_X5Y138_SLICE_X7Y138_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A6 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B1 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B2 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B4 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B5 = CLBLM_R_X5Y138_SLICE_X7Y138_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B6 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C2 = CLBLM_R_X5Y137_SLICE_X6Y137_D5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A1 = CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C4 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A2 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A3 = CLBLM_R_X5Y131_SLICE_X6Y131_C5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B1 = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B2 = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B3 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B4 = CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D2 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B5 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D5 = CLBLM_R_X5Y141_SLICE_X6Y141_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C1 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C2 = CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C3 = CLBLM_R_X5Y131_SLICE_X6Y131_D5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C4 = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C5 = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C6 = CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A4 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A5 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A6 = CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A3 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B1 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B2 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B3 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B5 = CLBLM_R_X7Y141_SLICE_X9Y141_CQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D2 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D3 = CLBLM_R_X3Y133_SLICE_X2Y133_B5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D4 = CLBLM_R_X3Y132_SLICE_X3Y132_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A1 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A2 = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C2 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A5 = CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C4 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C6 = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C3 = CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D1 = CLBLM_R_X5Y130_SLICE_X6Y130_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X13Y139_SLICE_X18Y139_BO5;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A1 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A2 = CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A3 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A6 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B1 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B2 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B4 = CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A1 = CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A2 = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A3 = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A5 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A6 = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C1 = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C2 = CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C3 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B1 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B3 = CLBLM_R_X3Y139_SLICE_X3Y139_CQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B5 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D2 = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D5 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D6 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B6 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C1 = CLBLL_L_X4Y133_SLICE_X5Y133_C5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C2 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C3 = CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A2 = CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A4 = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A6 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C6 = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_AX = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B1 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B4 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B6 = CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D2 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D4 = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D5 = CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C1 = CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C2 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C4 = CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C5 = CLBLM_L_X10Y140_SLICE_X12Y140_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C6 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A3 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A5 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A6 = CLBLL_L_X4Y131_SLICE_X4Y131_C5Q;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B1 = CLBLL_L_X2Y139_SLICE_X1Y139_CQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B2 = CLBLM_R_X3Y132_SLICE_X3Y132_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C2 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C3 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C4 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C5 = CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D1 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D2 = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D3 = CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D4 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D5 = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C1 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C5 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C6 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D3 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D5 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign LIOB33_X0Y63_IOB_X0Y64_O = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D6 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign RIOB33_X105Y151_IOB_X1Y152_O = 1'b1;
  assign RIOB33_X105Y151_IOB_X1Y151_O = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A6 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A1 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A5 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A6 = 1'b1;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C4 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A3 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A4 = CLBLM_R_X3Y134_SLICE_X3Y134_DQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A6 = CLBLM_R_X3Y135_SLICE_X2Y135_AO5;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C3 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B1 = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B2 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B4 = CLBLM_R_X3Y134_SLICE_X2Y134_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D1 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C4 = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C5 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D4 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D5 = CLBLL_L_X4Y133_SLICE_X4Y133_D5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A1 = CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A2 = CLBLM_R_X3Y134_SLICE_X3Y134_DQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A3 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A5 = CLBLM_R_X5Y134_SLICE_X7Y134_C5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_AX = CLBLM_R_X3Y135_SLICE_X2Y135_AO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B1 = CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B2 = CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B3 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B4 = CLBLM_R_X3Y134_SLICE_X3Y134_DQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B5 = CLBLM_R_X5Y131_SLICE_X6Y131_C5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C1 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C2 = CLBLM_R_X3Y134_SLICE_X2Y134_CQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C3 = CLBLL_L_X4Y133_SLICE_X4Y133_D5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C5 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C6 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D6 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B5 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C5 = CLBLM_R_X11Y141_SLICE_X14Y141_BO5;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C6 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D1 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D2 = CLBLM_R_X3Y134_SLICE_X2Y134_CQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D3 = CLBLM_R_X3Y134_SLICE_X2Y134_DQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D5 = CLBLL_L_X4Y131_SLICE_X4Y131_C5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A2 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A3 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A4 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B2 = CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y65_IOB_X0Y66_O = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A6 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign LIOB33_X0Y65_IOB_X0Y65_O = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign LIOB33_X0Y111_IOB_X0Y111_O = CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  assign RIOB33_X105Y153_IOB_X1Y154_O = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y153_O = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C2 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C3 = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C4 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C5 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C6 = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y159_IOB_X0Y160_O = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B4 = CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  assign LIOB33_X0Y159_IOB_X0Y159_O = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A1 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A2 = CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A3 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A5 = CLBLL_L_X2Y135_SLICE_X1Y135_BQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A6 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B2 = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B3 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B4 = CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B6 = CLBLL_L_X2Y135_SLICE_X1Y135_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B5 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C1 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C2 = CLBLM_R_X3Y134_SLICE_X2Y134_CQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C3 = CLBLM_R_X3Y134_SLICE_X2Y134_A5Q;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C4 = CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D2 = CLBLM_R_X3Y134_SLICE_X3Y134_DQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D3 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D5 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D6 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A1 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A3 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A4 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A5 = CLBLL_L_X2Y139_SLICE_X0Y139_B5Q;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_AX = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B1 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B2 = CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B3 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B4 = CLBLL_L_X2Y135_SLICE_X1Y135_DQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B5 = CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_BX = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C1 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C2 = CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C3 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C4 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C5 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C6 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D2 = CLBLM_R_X5Y144_SLICE_X7Y144_A5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_BX = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_C5Q;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C1 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign RIOB33_X105Y155_IOB_X1Y155_O = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D5 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C2 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D6 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign LIOB33_X0Y187_IOB_X0Y188_O = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign LIOB33_X0Y187_IOB_X0Y187_O = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C3 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C4 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C5 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D5 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B2 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D6 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A1 = CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A2 = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A3 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A5 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C6 = CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B3 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C1 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C2 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C4 = CLBLL_L_X2Y139_SLICE_X1Y139_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D2 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D4 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D5 = CLBLM_R_X3Y133_SLICE_X2Y133_CQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A1 = CLBLM_R_X3Y135_SLICE_X2Y135_BO5;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A3 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A4 = CLBLM_R_X3Y136_SLICE_X2Y136_DO5;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A6 = CLBLM_R_X7Y131_SLICE_X8Y131_BQ;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B1 = CLBLM_R_X3Y138_SLICE_X3Y138_DQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B2 = CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B4 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B5 = CLBLM_R_X3Y135_SLICE_X2Y135_AO5;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B6 = CLBLM_R_X3Y134_SLICE_X3Y134_DQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C1 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C2 = CLBLM_R_X3Y134_SLICE_X3Y134_DQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C3 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C4 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C5 = CLBLM_R_X3Y137_SLICE_X2Y137_DQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D1 = CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D2 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D3 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D4 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D5 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B6 = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C6 = CLBLM_R_X7Y133_SLICE_X8Y133_DO5;
  assign RIOB33_X105Y157_IOB_X1Y157_O = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y158_O = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y189_IOB_X0Y190_O = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign LIOB33_X0Y189_IOB_X0Y189_O = CLBLL_L_X2Y139_SLICE_X0Y139_AQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D5 = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A3 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A5 = CLBLM_R_X3Y134_SLICE_X3Y134_D5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A6 = CLBLL_L_X2Y139_SLICE_X1Y139_DQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B2 = CLBLM_R_X3Y137_SLICE_X3Y137_DQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B4 = CLBLM_R_X7Y137_SLICE_X8Y137_B5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B5 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C2 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C3 = CLBLM_R_X5Y141_SLICE_X6Y141_B5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C5 = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D1 = CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D3 = CLBLL_L_X2Y137_SLICE_X1Y137_C5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D4 = CLBLM_R_X3Y135_SLICE_X3Y135_C5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D5 = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A1 = CLBLM_R_X3Y135_SLICE_X2Y135_BO5;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A3 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A4 = CLBLM_R_X3Y136_SLICE_X2Y136_DO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A5 = CLBLL_L_X4Y138_SLICE_X5Y138_CQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A6 = CLBLM_R_X3Y134_SLICE_X3Y134_DQ;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B1 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B2 = CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B3 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B4 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B6 = CLBLM_R_X3Y137_SLICE_X3Y137_B5Q;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C2 = CLBLM_R_X3Y137_SLICE_X2Y137_CQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C3 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C4 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C6 = CLBLL_L_X4Y135_SLICE_X5Y135_A5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D1 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D3 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D4 = CLBLM_R_X3Y138_SLICE_X2Y138_A5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOB33_X105Y159_IOB_X1Y160_O = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y159_O = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D6 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y192_O = CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  assign LIOB33_X0Y191_IOB_X0Y191_O = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_R_X5Y138_SLICE_X7Y138_A5Q;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A1 = CLBLM_R_X3Y136_SLICE_X3Y136_B5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A3 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A4 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A5 = CLBLM_R_X5Y137_SLICE_X6Y137_B5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B1 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B2 = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B4 = CLBLL_L_X2Y139_SLICE_X0Y139_BQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B5 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C1 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C3 = CLBLM_R_X3Y138_SLICE_X3Y138_D5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C4 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C5 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D1 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D2 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D4 = CLBLL_L_X4Y137_SLICE_X4Y137_C5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A1 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A3 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A5 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B1 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B2 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B3 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B4 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C1 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C2 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C3 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C5 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C6 = CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D2 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D3 = CLBLM_R_X3Y138_SLICE_X2Y138_DQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D6 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_R_X5Y138_SLICE_X7Y138_A5Q;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y194_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOB33_X0Y193_IOB_X0Y193_O = CLBLM_R_X3Y165_SLICE_X2Y165_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C3 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A2 = CLBLM_R_X3Y139_SLICE_X3Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A3 = CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A6 = CLBLM_R_X3Y138_SLICE_X2Y138_A5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C4 = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_AX = CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B2 = CLBLM_R_X3Y138_SLICE_X3Y138_DQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B3 = CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B4 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C6 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C1 = CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C3 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C4 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C5 = CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D1 = CLBLM_R_X3Y139_SLICE_X3Y139_C5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D2 = CLBLL_L_X2Y139_SLICE_X1Y139_DQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D3 = CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D4 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D5 = CLBLM_R_X3Y139_SLICE_X2Y139_CO5;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D6 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A2 = CLBLM_R_X3Y139_SLICE_X3Y139_B5Q;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A3 = CLBLM_R_X3Y140_SLICE_X2Y140_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A4 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A5 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_AX = CLBLM_R_X3Y140_SLICE_X2Y140_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B1 = CLBLL_L_X2Y139_SLICE_X1Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B2 = CLBLL_L_X2Y139_SLICE_X1Y139_CQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B3 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B4 = CLBLL_L_X2Y139_SLICE_X1Y139_DQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B5 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D2 = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C1 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C2 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C3 = CLBLL_L_X2Y139_SLICE_X1Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C5 = CLBLL_L_X2Y139_SLICE_X1Y139_CQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_R_X5Y138_SLICE_X7Y138_B5Q;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D2 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D3 = CLBLM_R_X3Y137_SLICE_X3Y137_B5Q;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D4 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D5 = CLBLM_R_X3Y139_SLICE_X3Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D6 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D4 = CLBLM_R_X11Y136_SLICE_X14Y136_AO5;
  assign LIOB33_X0Y195_IOB_X0Y195_O = CLBLM_R_X3Y140_SLICE_X2Y140_CO5;
  assign LIOB33_X0Y195_IOB_X0Y196_O = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D5 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A1 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A3 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A4 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A6 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B6 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y162_O = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C6 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y161_O = CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A5 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C5 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C6 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A1 = CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A2 = CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A3 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A5 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A6 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B1 = CLBLM_R_X3Y140_SLICE_X3Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B2 = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B3 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B5 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B6 = CLBLM_R_X3Y138_SLICE_X3Y138_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C1 = CLBLM_R_X3Y137_SLICE_X3Y137_C5Q;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C2 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C4 = CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C5 = CLBLM_R_X3Y140_SLICE_X3Y140_DO5;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D6 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_C5Q;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D3 = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D4 = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D5 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = CLBLM_R_X13Y139_SLICE_X18Y139_AO6;
  assign RIOB33_X105Y165_IOB_X1Y166_O = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A2 = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A3 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A4 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A6 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_AX = CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B2 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B3 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B4 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B5 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B6 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C1 = CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C2 = CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C3 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C4 = CLBLM_R_X3Y135_SLICE_X2Y135_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D1 = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D3 = CLBLM_R_X3Y136_SLICE_X3Y136_B5Q;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D4 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D6 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y197_O = CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B6 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A1 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A2 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A3 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A5 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B1 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B3 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B5 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A2 = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A3 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A4 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A5 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y167_O = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B2 = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B3 = CLBLM_R_X3Y138_SLICE_X3Y138_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B4 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B5 = CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B6 = CLBLL_L_X4Y141_SLICE_X4Y141_DQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C1 = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C2 = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C3 = CLBLL_L_X4Y140_SLICE_X4Y140_C5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C4 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C5 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C6 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D2 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D3 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D4 = CLBLL_L_X4Y140_SLICE_X4Y140_C5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D5 = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D6 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A1 = CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A2 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A3 = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A4 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A6 = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B1 = CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B2 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B3 = CLBLL_L_X4Y141_SLICE_X4Y141_DQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B4 = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B6 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C3 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C6 = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C4 = CLBLM_L_X10Y140_SLICE_X12Y140_DO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A2 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A3 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A4 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A5 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B2 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B3 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B4 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B5 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C2 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C3 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C4 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C5 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D2 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D3 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D4 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D5 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A3 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A5 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B2 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B5 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B6 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C2 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C3 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C4 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C5 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D2 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D3 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D4 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D5 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D6 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A2 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A3 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A4 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A5 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A6 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A2 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A4 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A2 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A4 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B2 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C1 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C2 = CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C3 = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C4 = CLBLM_R_X5Y133_SLICE_X6Y133_DQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C5 = CLBLM_L_X12Y137_SLICE_X16Y137_BO5;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C6 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D1 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D3 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D6 = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_A5Q;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X4Y131_SLICE_X5Y131_D5Q;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B3 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B4 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B5 = CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B6 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C6 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A1 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A2 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A3 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A4 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A5 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A6 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B1 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B2 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B3 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B4 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B5 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B6 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C1 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C2 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C3 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C4 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C5 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D1 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D2 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D3 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D4 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D5 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D6 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A2 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A3 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A5 = CLBLM_R_X7Y139_SLICE_X8Y139_CQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A6 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B2 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B3 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B6 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C2 = CLBLM_R_X11Y138_SLICE_X14Y138_AO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C3 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C4 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C5 = CLBLM_L_X12Y138_SLICE_X16Y138_BO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C6 = CLBLM_R_X11Y139_SLICE_X14Y139_DO5;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D1 = CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D2 = CLBLM_R_X7Y139_SLICE_X8Y139_CQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D5 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D6 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C6 = CLBLM_L_X10Y134_SLICE_X13Y134_C5Q;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A2 = CLBLM_L_X10Y138_SLICE_X12Y138_CQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A4 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B2 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B6 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D1 = CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C2 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C6 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D2 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D6 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A1 = CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A2 = CLBLM_L_X10Y138_SLICE_X12Y138_CQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A5 = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A6 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B2 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B6 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C2 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D2 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_D1 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_D1 = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A1 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A3 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A4 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A5 = CLBLM_L_X10Y134_SLICE_X13Y134_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A6 = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C6 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLL_L_X2Y139_SLICE_X0Y139_AQ;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D6 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = CLBLM_R_X13Y139_SLICE_X18Y139_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A1 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A2 = CLBLM_R_X7Y133_SLICE_X9Y133_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A6 = CLBLM_R_X11Y134_SLICE_X14Y134_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B3 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B4 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B5 = CLBLM_L_X8Y139_SLICE_X10Y139_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B6 = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C2 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C4 = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D3 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D6 = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = CLBLL_L_X2Y139_SLICE_X0Y139_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A1 = CLBLM_L_X8Y139_SLICE_X11Y139_DQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A3 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A4 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A6 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B1 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B2 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B4 = CLBLM_R_X5Y138_SLICE_X7Y138_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B5 = CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B6 = CLBLM_L_X10Y133_SLICE_X12Y133_A5Q;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C1 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C2 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C3 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D1 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D2 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D4 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D5 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D6 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A1 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A3 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A6 = CLBLM_L_X10Y133_SLICE_X12Y133_A5Q;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_R_X5Y138_SLICE_X7Y138_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B1 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B2 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B3 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B5 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B6 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C1 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C2 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C6 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D1 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D2 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D5 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D6 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B2 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B3 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B5 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B6 = CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C2 = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign RIOB33_X105Y183_IOB_X1Y183_O = 1'b0;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A2 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A3 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A4 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A6 = CLBLM_R_X3Y129_SLICE_X3Y129_BO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B2 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B3 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B4 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B6 = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C1 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C2 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C3 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C4 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C5 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A3 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A4 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_C5Q;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D1 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D2 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D3 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D4 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D5 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D6 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A6 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B1 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B3 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B4 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B6 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C1 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C2 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C4 = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C5 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C6 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D1 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D2 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D5 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D6 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A1 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A2 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A3 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A4 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A6 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A1 = CLBLM_L_X10Y134_SLICE_X12Y134_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A3 = CLBLM_R_X3Y134_SLICE_X3Y134_C5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A5 = CLBLM_R_X5Y138_SLICE_X7Y138_A5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B2 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B3 = CLBLL_L_X4Y129_SLICE_X4Y129_CO5;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B4 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C2 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C4 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C5 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C6 = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B1 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B4 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B5 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B6 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C1 = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D3 = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D5 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C4 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C5 = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D1 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D2 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D3 = CLBLM_L_X10Y134_SLICE_X12Y134_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D5 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D6 = CLBLM_L_X8Y140_SLICE_X10Y140_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D4 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X13Y139_SLICE_X18Y139_AO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A5 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A6 = CLBLL_L_X4Y141_SLICE_X4Y141_CQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A2 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A3 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A5 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A6 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B1 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B2 = CLBLM_L_X10Y134_SLICE_X13Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B3 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B5 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C1 = CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C2 = CLBLM_L_X10Y134_SLICE_X13Y134_CQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C3 = CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C5 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D1 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D2 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D3 = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D4 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D5 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D6 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A2 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A3 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A4 = CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A6 = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B1 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B2 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B3 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C2 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C3 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C4 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C5 = CLBLM_L_X10Y137_SLICE_X12Y137_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C6 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D1 = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D2 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D3 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D4 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D5 = CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D6 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLM_R_X5Y130_SLICE_X6Y130_CQ;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A3 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A4 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A6 = CLBLM_R_X3Y133_SLICE_X2Y133_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_AX = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B3 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B5 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_BX = CLBLL_L_X4Y131_SLICE_X4Y131_DO5;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C1 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C2 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C5 = CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D1 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D2 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D5 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A2 = CLBLM_R_X7Y137_SLICE_X9Y137_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A4 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A5 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B2 = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B4 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B5 = CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C2 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C3 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C5 = CLBLM_R_X7Y137_SLICE_X9Y137_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C6 = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A2 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A3 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D1 = CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D2 = CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D3 = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D4 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D5 = CLBLM_L_X10Y135_SLICE_X12Y135_DQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D6 = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A5 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A6 = CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B2 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B3 = CLBLL_L_X4Y136_SLICE_X4Y136_C5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B4 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B5 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B6 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C2 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C4 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B2 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B3 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B4 = CLBLM_R_X11Y134_SLICE_X14Y134_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B5 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B6 = CLBLM_R_X3Y136_SLICE_X3Y136_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D2 = CLBLL_L_X4Y133_SLICE_X5Y133_C5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C1 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C4 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D5 = CLBLM_R_X5Y133_SLICE_X7Y133_B5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D2 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D3 = CLBLM_L_X10Y135_SLICE_X12Y135_DQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D4 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D6 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A3 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A6 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B3 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B6 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLM_R_X3Y139_SLICE_X3Y139_CQ;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C3 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C6 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D3 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D6 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A3 = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_CQ;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A6 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X13Y139_SLICE_X18Y139_AO5;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B3 = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B4 = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B5 = CLBLM_L_X10Y138_SLICE_X12Y138_CQ;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B6 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_CQ;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C3 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C4 = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C6 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D3 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A1 = CLBLL_L_X4Y133_SLICE_X4Y133_DQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A3 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B1 = CLBLL_L_X4Y136_SLICE_X4Y136_B5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B4 = CLBLM_R_X5Y132_SLICE_X6Y132_A5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B6 = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C2 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C3 = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C5 = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D3 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A1 = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A2 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_D5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A4 = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A5 = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A6 = CLBLM_R_X3Y137_SLICE_X2Y137_CQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_AX = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B1 = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B2 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B3 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B4 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B5 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B6 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C1 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C2 = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C3 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C4 = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C5 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C6 = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A1 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A2 = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A3 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A5 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A6 = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B1 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B2 = CLBLL_L_X4Y133_SLICE_X4Y133_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B5 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B6 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D1 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D2 = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D3 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C1 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C2 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A1 = CLBLM_L_X10Y137_SLICE_X12Y137_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C3 = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C4 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C5 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C6 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A3 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A4 = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B1 = CLBLM_R_X5Y142_SLICE_X7Y142_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D2 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D3 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D4 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D5 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D6 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B2 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C1 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C2 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B5 = CLBLM_L_X10Y139_SLICE_X13Y139_DQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B6 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C3 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D2 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D3 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D4 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D5 = CLBLM_L_X10Y138_SLICE_X12Y138_B5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D6 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_R_X13Y139_SLICE_X18Y139_CO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = CLBLM_R_X3Y140_SLICE_X2Y140_CO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X2Y137_SLICE_X0Y137_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A1 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A2 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A3 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A5 = CLBLL_L_X4Y139_SLICE_X4Y139_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A6 = CLBLM_R_X3Y133_SLICE_X2Y133_C5Q;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B1 = CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B2 = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B3 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C1 = CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C3 = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C5 = CLBLL_L_X4Y133_SLICE_X4Y133_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D1 = CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D2 = CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D3 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A1 = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A2 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A3 = CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A4 = CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A5 = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B1 = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B2 = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B3 = CLBLM_L_X10Y134_SLICE_X13Y134_C5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B4 = CLBLM_R_X7Y140_SLICE_X8Y140_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B5 = CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B6 = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A1 = CLBLL_L_X4Y133_SLICE_X5Y133_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C3 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C4 = CLBLM_R_X7Y140_SLICE_X8Y140_CQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A3 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A4 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A5 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C5 = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B2 = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B4 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B5 = CLBLL_L_X4Y141_SLICE_X4Y141_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D3 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D4 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C1 = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C2 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C4 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C5 = CLBLM_R_X7Y132_SLICE_X8Y132_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D6 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A5 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A2 = CLBLL_L_X4Y138_SLICE_X5Y138_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D2 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B1 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B3 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B4 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B5 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D3 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D4 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C1 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C3 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C4 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C5 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLM_R_X3Y132_SLICE_X3Y132_A5Q;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X4Y131_SLICE_X5Y131_D5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D1 = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D2 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D3 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D5 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D6 = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X13Y139_SLICE_X18Y139_CO6;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A1 = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A2 = CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A4 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B1 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B3 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B4 = CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C1 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C2 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C3 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C4 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C5 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D1 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D2 = CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D3 = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D4 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D5 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D6 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A1 = CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A2 = CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A3 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A4 = CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A5 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A6 = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_AX = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B4 = CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B6 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A2 = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A3 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C1 = CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C2 = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C3 = CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C4 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C5 = CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C6 = CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A4 = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B1 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B2 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D1 = CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D2 = CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D3 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D4 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D5 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D6 = CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C1 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C2 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C3 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C4 = CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C5 = CLBLL_L_X4Y134_SLICE_X5Y134_BO5;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A1 = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A2 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D3 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D4 = CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D5 = CLBLL_L_X4Y134_SLICE_X5Y134_BO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D6 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B1 = CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B4 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C1 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C2 = CLBLM_R_X3Y138_SLICE_X2Y138_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C3 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C4 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D2 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_DQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D5 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D6 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A1 = CLBLL_L_X4Y133_SLICE_X4Y133_DQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A2 = CLBLM_R_X5Y140_SLICE_X6Y140_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A3 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A4 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B1 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B3 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B4 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B5 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C2 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C3 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C4 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C5 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C6 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D2 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D3 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D4 = CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D5 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A1 = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A2 = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A4 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A5 = CLBLM_R_X3Y133_SLICE_X2Y133_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B1 = CLBLM_L_X8Y139_SLICE_X11Y139_DQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B2 = CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A1 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A2 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B4 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B5 = CLBLM_L_X10Y138_SLICE_X12Y138_CQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B6 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A3 = CLBLM_R_X5Y130_SLICE_X6Y130_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_BX = CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A5 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C2 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C3 = CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C4 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B1 = CLBLM_R_X3Y137_SLICE_X2Y137_DQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C1 = CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B4 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C4 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D3 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D4 = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D5 = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C3 = CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C5 = CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_D5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D2 = CLBLL_L_X2Y138_SLICE_X1Y138_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D3 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D4 = CLBLM_R_X5Y133_SLICE_X7Y133_B5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D5 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D6 = CLBLL_L_X2Y138_SLICE_X1Y138_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A1 = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_AX = CLBLM_R_X3Y137_SLICE_X2Y137_CQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A3 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B1 = CLBLM_L_X10Y139_SLICE_X13Y139_DQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X11Y139_SLICE_X14Y139_CO5;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_BX = CLBLM_R_X5Y139_SLICE_X6Y139_CQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C3 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D1 = CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D2 = CLBLM_L_X8Y132_SLICE_X10Y132_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D3 = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D4 = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D5 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D6 = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A5 = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A1 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A2 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A5 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A6 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C6 = 1'b1;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D6 = 1'b1;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A2 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A3 = CLBLL_L_X4Y140_SLICE_X5Y140_C5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A5 = CLBLM_R_X3Y136_SLICE_X3Y136_D5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B3 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B4 = CLBLM_L_X8Y140_SLICE_X10Y140_B5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B5 = CLBLL_L_X4Y136_SLICE_X4Y136_C5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C1 = CLBLM_R_X5Y141_SLICE_X6Y141_C5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C3 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C4 = CLBLL_L_X4Y131_SLICE_X5Y131_D5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C5 = CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D1 = CLBLL_L_X2Y138_SLICE_X1Y138_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D2 = CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_B5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D5 = CLBLL_L_X4Y135_SLICE_X4Y135_B5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign LIOB33_X0Y113_IOB_X0Y113_O = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A1 = CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A3 = CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A4 = CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A5 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A1 = CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A3 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A4 = CLBLM_R_X3Y134_SLICE_X2Y134_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A6 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_AX = CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B1 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B2 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B2 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B4 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B5 = CLBLL_L_X4Y140_SLICE_X5Y140_C5Q;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C2 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C3 = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C5 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A6 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B4 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D1 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D2 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D3 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D6 = CLBLM_R_X3Y140_SLICE_X2Y140_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B1 = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B2 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A2 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A5 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A6 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_BX = CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C2 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C3 = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B2 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B3 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B5 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B6 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_CX = CLBLM_R_X11Y140_SLICE_X14Y140_AO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D2 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C1 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C2 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C3 = CLBLM_L_X8Y131_SLICE_X10Y131_D5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C5 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C6 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D4 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D2 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D3 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D4 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D6 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A2 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A4 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A5 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B5 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B6 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C1 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C2 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C3 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C4 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C5 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C6 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D1 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D2 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D4 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D5 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D6 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A3 = CLBLM_R_X7Y138_SLICE_X8Y138_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A4 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B1 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B3 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C1 = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C3 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C4 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C6 = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D1 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D2 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D3 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D4 = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D6 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A1 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A3 = CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A4 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A5 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B1 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B2 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B3 = CLBLM_L_X10Y135_SLICE_X12Y135_DQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B4 = CLBLM_R_X3Y138_SLICE_X2Y138_BQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B6 = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C1 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C3 = CLBLM_R_X3Y137_SLICE_X2Y137_D5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C4 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C5 = CLBLL_L_X4Y141_SLICE_X4Y141_DQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C6 = 1'b1;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X5Y138_SLICE_X6Y138_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D1 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D2 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D3 = CLBLL_L_X4Y136_SLICE_X5Y136_DQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A1 = CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A1 = CLBLM_R_X3Y133_SLICE_X2Y133_B5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A2 = CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A3 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A4 = CLBLL_L_X4Y137_SLICE_X5Y137_DQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A5 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A2 = CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A3 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B1 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B1 = CLBLM_R_X5Y140_SLICE_X6Y140_B5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B2 = CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B3 = CLBLL_L_X4Y137_SLICE_X5Y137_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B4 = CLBLL_L_X4Y137_SLICE_X5Y137_DQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B5 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B3 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A2 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A3 = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A4 = CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A5 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C2 = CLBLM_R_X5Y140_SLICE_X7Y140_D5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C3 = CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C4 = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A6 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C5 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B4 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B2 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B3 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B6 = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D1 = CLBLM_R_X5Y141_SLICE_X6Y141_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D3 = CLBLL_L_X4Y137_SLICE_X5Y137_DQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D4 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D5 = CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C1 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C4 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C5 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D1 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D2 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D3 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D4 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D5 = CLBLM_R_X5Y133_SLICE_X7Y133_B5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D6 = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A6 = CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B2 = CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B3 = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A4 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A6 = CLBLM_R_X7Y133_SLICE_X9Y133_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C1 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C2 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B2 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B4 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B5 = CLBLM_R_X5Y135_SLICE_X7Y135_B5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D1 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D2 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C1 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C2 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C4 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C5 = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D3 = CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D5 = CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D6 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D3 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D4 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D5 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y138_SLICE_X5Y138_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X2Y139_SLICE_X0Y139_BQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A1 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A2 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A4 = CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A5 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A6 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = CLBLM_R_X3Y133_SLICE_X2Y133_DO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B1 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B2 = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B3 = CLBLM_L_X10Y134_SLICE_X13Y134_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B4 = CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B5 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B6 = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C1 = CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C2 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C3 = CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C4 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C5 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C6 = CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D1 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D2 = CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D3 = CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D4 = CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D5 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D6 = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A1 = CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A2 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A3 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A5 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B5 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B1 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B6 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B2 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B4 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B5 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C1 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C2 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C3 = CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C4 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C5 = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C6 = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D1 = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D2 = CLBLM_R_X7Y141_SLICE_X9Y141_C5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D3 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C1 = CLBLM_R_X5Y137_SLICE_X6Y137_C5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D5 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D6 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A1 = CLBLM_R_X3Y138_SLICE_X3Y138_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A2 = CLBLL_L_X2Y139_SLICE_X0Y139_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A3 = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A4 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A5 = CLBLM_R_X5Y137_SLICE_X6Y137_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A6 = CLBLL_L_X4Y138_SLICE_X5Y138_CQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_AX = CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B1 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B2 = CLBLM_R_X5Y135_SLICE_X7Y135_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B3 = CLBLM_R_X3Y138_SLICE_X3Y138_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B4 = CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B5 = CLBLL_L_X4Y137_SLICE_X4Y137_C5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B6 = CLBLM_R_X5Y134_SLICE_X7Y134_DQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C1 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C2 = CLBLM_R_X7Y137_SLICE_X8Y137_C5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C3 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C5 = CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C6 = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D2 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D3 = CLBLM_R_X3Y138_SLICE_X3Y138_CQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D5 = CLBLM_R_X7Y138_SLICE_X8Y138_A5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D6 = CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A2 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A3 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A5 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A1 = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A3 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B1 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B2 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B4 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A5 = CLBLM_L_X10Y134_SLICE_X13Y134_C5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C1 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C2 = CLBLM_R_X3Y138_SLICE_X3Y138_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C3 = CLBLM_L_X10Y138_SLICE_X12Y138_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C4 = CLBLL_L_X4Y140_SLICE_X5Y140_A5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A1 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A2 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A5 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A3 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B1 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B3 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B4 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B5 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D6 = CLBLL_L_X2Y138_SLICE_X1Y138_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D1 = CLBLL_L_X2Y138_SLICE_X1Y138_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C1 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C2 = CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C3 = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C5 = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C4 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D4 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A2 = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A3 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A4 = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A5 = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D2 = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D3 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D5 = CLBLM_L_X8Y131_SLICE_X11Y131_C5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D6 = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B1 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B2 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B3 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A2 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A4 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C1 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C2 = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B1 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B2 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B3 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B5 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C1 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C2 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C3 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C4 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D2 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D3 = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D4 = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D5 = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A1 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A2 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A3 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A4 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A5 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B1 = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B2 = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B3 = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B4 = CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B5 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B6 = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C1 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C2 = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C3 = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C4 = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C6 = CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D1 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D2 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D3 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D4 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D5 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D6 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A1 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A3 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A5 = CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B1 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B4 = CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B5 = CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B6 = CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X13Y139_SLICE_X18Y139_BO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C1 = CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C2 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C3 = CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C4 = CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C5 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C6 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D1 = CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D2 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D3 = CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D4 = CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A1 = CLBLM_R_X5Y141_SLICE_X6Y141_B5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A2 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A3 = CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A4 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D5 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D6 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B1 = CLBLL_L_X4Y140_SLICE_X4Y140_DQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B3 = CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B4 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B5 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B6 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C1 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C3 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C5 = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C6 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D1 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D2 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D3 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D4 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D5 = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D6 = CLBLM_R_X5Y132_SLICE_X6Y132_A5Q;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A1 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A2 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A3 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A4 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A5 = CLBLL_L_X4Y137_SLICE_X5Y137_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C2 = CLBLL_L_X4Y140_SLICE_X4Y140_C5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A1 = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B1 = CLBLL_L_X4Y139_SLICE_X5Y139_CQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B2 = CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B3 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A5 = CLBLM_R_X5Y144_SLICE_X7Y144_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A6 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B4 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B5 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A2 = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A3 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B2 = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B3 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B6 = CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C1 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C2 = CLBLL_L_X4Y139_SLICE_X5Y139_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C1 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C2 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C3 = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C4 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C5 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C6 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A1 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A3 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D2 = CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D3 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D5 = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D6 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C1 = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C2 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C3 = CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C4 = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C6 = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C5 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A2 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A3 = CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A5 = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D1 = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D2 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D3 = CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D4 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D5 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B5 = CLBLM_R_X5Y140_SLICE_X7Y140_C5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B6 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D6 = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B1 = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B2 = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B3 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A1 = CLBLM_L_X8Y131_SLICE_X10Y131_DQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C4 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C5 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A2 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A3 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A4 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A6 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B1 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B2 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B5 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D2 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C1 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C2 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C3 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C4 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C6 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D5 = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D1 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D2 = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D3 = CLBLM_R_X3Y133_SLICE_X2Y133_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D4 = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D6 = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A1 = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A2 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A3 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A5 = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A6 = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B1 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B2 = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B3 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B4 = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B5 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B6 = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C1 = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C2 = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C3 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C4 = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C5 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C6 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D1 = CLBLM_L_X10Y137_SLICE_X13Y137_AO5;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D2 = CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D3 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D4 = CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D5 = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D6 = CLBLM_L_X10Y138_SLICE_X12Y138_C5Q;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A1 = CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A2 = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A3 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A5 = CLBLM_L_X8Y140_SLICE_X11Y140_C5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B1 = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B2 = CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B3 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B4 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B5 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B6 = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C1 = CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C3 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C4 = CLBLM_L_X10Y139_SLICE_X12Y139_AO5;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C5 = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C6 = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B3 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A2 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A3 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A4 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A6 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B4 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B5 = CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B1 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B2 = CLBLM_R_X5Y141_SLICE_X6Y141_C5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B3 = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B5 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C1 = CLBLL_L_X4Y140_SLICE_X4Y140_C5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C2 = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C4 = CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C5 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_BX = CLBLM_L_X8Y131_SLICE_X11Y131_C5Q;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D2 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D3 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D4 = CLBLM_R_X3Y138_SLICE_X2Y138_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D5 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D6 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C1 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C2 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C4 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C5 = CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = CLBLM_R_X3Y165_SLICE_X2Y165_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A1 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A2 = CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A4 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A5 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B1 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B2 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B4 = CLBLL_L_X4Y140_SLICE_X5Y140_CQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B5 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C1 = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C2 = CLBLM_R_X5Y139_SLICE_X6Y139_CQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C3 = CLBLM_R_X7Y140_SLICE_X8Y140_B5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C4 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A1 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A2 = CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A3 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A6 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D2 = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D4 = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B1 = CLBLM_R_X5Y135_SLICE_X6Y135_DQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D5 = CLBLM_R_X3Y135_SLICE_X3Y135_C5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B5 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B4 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B2 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C1 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C2 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C3 = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C4 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C5 = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C6 = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D3 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D2 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D3 = CLBLM_L_X10Y135_SLICE_X12Y135_C5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D5 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A1 = CLBLM_L_X8Y131_SLICE_X10Y131_DQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A2 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B1 = CLBLM_R_X7Y131_SLICE_X9Y131_B5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B2 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B3 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B5 = CLBLM_L_X10Y134_SLICE_X13Y134_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C1 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C3 = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C4 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C5 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C6 = CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A2 = CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D1 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D3 = CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D4 = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D5 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A3 = CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C6 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A5 = CLBLM_L_X8Y139_SLICE_X11Y139_D5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A2 = CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A3 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A5 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A6 = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B1 = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B2 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B3 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B5 = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B6 = CLBLM_R_X11Y138_SLICE_X15Y138_AO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B4 = CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C2 = CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C3 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C4 = CLBLM_R_X11Y138_SLICE_X15Y138_AO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B5 = CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C5 = CLBLM_R_X11Y138_SLICE_X14Y138_AO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C6 = CLBLM_L_X12Y138_SLICE_X16Y138_AO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B6 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D1 = CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D2 = CLBLM_R_X11Y139_SLICE_X15Y139_AO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_C5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D4 = CLBLM_R_X3Y139_SLICE_X3Y139_B5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D5 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A1 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A2 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A3 = CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A6 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B1 = CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B2 = CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B3 = CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B4 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B5 = CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C1 = CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C2 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C3 = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C4 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C5 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C6 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C4 = CLBLM_L_X8Y140_SLICE_X11Y140_C5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A2 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A3 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A4 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A6 = CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C5 = CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C6 = CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B1 = CLBLL_L_X4Y140_SLICE_X4Y140_DQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B2 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B3 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B4 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B5 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D2 = CLBLM_R_X11Y139_SLICE_X15Y139_BO5;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D3 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C1 = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C3 = CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C5 = CLBLL_L_X4Y140_SLICE_X5Y140_C5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B4 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D1 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D2 = CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D3 = CLBLL_L_X4Y141_SLICE_X4Y141_DQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D4 = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D5 = CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B5 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A2 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A3 = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A4 = CLBLL_L_X4Y136_SLICE_X5Y136_C5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B1 = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B2 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B3 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B4 = CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B5 = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B6 = CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C1 = CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C2 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C4 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C5 = CLBLM_R_X3Y139_SLICE_X3Y139_C5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D1 = CLBLM_R_X5Y140_SLICE_X7Y140_D5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D3 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D4 = CLBLM_R_X5Y138_SLICE_X6Y138_C5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D5 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A1 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A2 = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A4 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A5 = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A6 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B1 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B3 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B4 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B5 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B6 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C1 = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C2 = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C3 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C4 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C5 = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D1 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D2 = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D4 = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D5 = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D6 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A2 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A4 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D2 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B1 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B2 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B3 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B4 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B5 = CLBLL_L_X4Y133_SLICE_X4Y133_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C1 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C2 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C3 = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C5 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D2 = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_BO5;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D4 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D5 = CLBLM_R_X7Y131_SLICE_X9Y131_B5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D6 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A1 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A3 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A5 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B1 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B2 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B5 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A1 = CLBLM_L_X8Y131_SLICE_X10Y131_D5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A2 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A3 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C1 = CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C3 = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D1 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D2 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D3 = CLBLM_R_X3Y139_SLICE_X3Y139_B5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A2 = CLBLM_L_X10Y139_SLICE_X12Y139_AO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A3 = CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A4 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A6 = CLBLM_L_X10Y139_SLICE_X12Y139_BO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B1 = CLBLM_L_X10Y139_SLICE_X13Y139_DQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B4 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A1 = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A2 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A3 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A6 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_AX = CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B1 = CLBLM_R_X7Y141_SLICE_X9Y141_CQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B2 = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B3 = CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B4 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B5 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C1 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C3 = CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C4 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C5 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A3 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D3 = CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D4 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D6 = CLBLM_R_X3Y139_SLICE_X3Y139_C5Q;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_R_X13Y139_SLICE_X18Y139_CO5;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A1 = CLBLM_R_X5Y142_SLICE_X7Y142_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A3 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A4 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A5 = CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A6 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B2 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B4 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B6 = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C1 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C2 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C3 = CLBLM_R_X3Y139_SLICE_X3Y139_C5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C4 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C5 = CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C6 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D4 = CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D5 = CLBLL_L_X4Y136_SLICE_X5Y136_C5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D6 = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A2 = CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A3 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A5 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B4 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B6 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C1 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C2 = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C3 = CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C4 = CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D1 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D2 = CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D3 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D4 = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D5 = CLBLM_L_X8Y138_SLICE_X11Y138_BO5;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A1 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A2 = CLBLM_L_X8Y139_SLICE_X11Y139_DQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A3 = CLBLM_L_X8Y134_SLICE_X11Y134_DO5;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A4 = CLBLM_R_X5Y141_SLICE_X6Y141_DO5;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A5 = CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A6 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_AX = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B1 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B2 = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B4 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B5 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C1 = CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C2 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C3 = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C4 = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C5 = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C6 = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D1 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D2 = CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D3 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D4 = CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D5 = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D6 = CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A2 = CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A3 = CLBLM_R_X5Y135_SLICE_X7Y135_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A4 = CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A5 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B1 = CLBLM_L_X12Y138_SLICE_X16Y138_DO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B2 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B3 = CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B4 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B6 = CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A2 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A3 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A5 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A6 = CLBLM_R_X3Y140_SLICE_X3Y140_A5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B3 = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B5 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C1 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C2 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C3 = CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C5 = CLBLM_R_X5Y142_SLICE_X7Y142_D5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D3 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A2 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A3 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A4 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B6 = CLBLM_L_X10Y139_SLICE_X12Y139_BO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A5 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_AX = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B2 = CLBLM_R_X7Y141_SLICE_X9Y141_C5Q;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B3 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A3 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A4 = CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A5 = CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A6 = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A1 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A2 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A3 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B2 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B3 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B4 = CLBLM_R_X7Y130_SLICE_X8Y130_DO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B5 = CLBLM_R_X3Y134_SLICE_X3Y134_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B6 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_AX = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B1 = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C1 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C2 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C4 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C5 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C6 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_BX = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C1 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C3 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C4 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C6 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D3 = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D4 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D5 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D6 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D6 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A1 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A2 = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A3 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A4 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A5 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B1 = CLBLL_L_X4Y141_SLICE_X4Y141_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B2 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B5 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C1 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C2 = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C3 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C4 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C5 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D3 = CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D4 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D6 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A1 = CLBLM_R_X7Y133_SLICE_X9Y133_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A3 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A6 = CLBLM_L_X10Y138_SLICE_X12Y138_C5Q;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B2 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B3 = CLBLM_L_X8Y134_SLICE_X10Y134_B5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B4 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B5 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B6 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_CQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C1 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C2 = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C3 = CLBLM_R_X7Y137_SLICE_X8Y137_B5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C4 = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C5 = CLBLM_R_X5Y137_SLICE_X6Y137_D5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C6 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D1 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D2 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D3 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D4 = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D5 = CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D6 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C2 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A2 = CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A3 = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A4 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A5 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A6 = CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B1 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B2 = CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B3 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B4 = CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B6 = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C3 = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C1 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C2 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C3 = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C4 = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C5 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C6 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D1 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D3 = CLBLM_R_X7Y134_SLICE_X8Y134_DQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D4 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C4 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A1 = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A2 = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A3 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A4 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A6 = CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B2 = CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B3 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B4 = CLBLM_R_X11Y141_SLICE_X14Y141_BO5;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B5 = CLBLM_L_X10Y140_SLICE_X13Y140_BO5;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B6 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A1 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A3 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A4 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C4 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B3 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B4 = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B5 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D1 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C1 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C2 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C4 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D2 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D4 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A1 = CLBLM_R_X7Y134_SLICE_X8Y134_DQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A2 = CLBLM_L_X10Y140_SLICE_X13Y140_BO5;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D3 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A3 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A4 = CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D1 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D4 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D3 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D4 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D6 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D2 = CLBLM_R_X7Y131_SLICE_X8Y131_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D5 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B1 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B2 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B3 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A2 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A3 = CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A4 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A6 = CLBLL_L_X4Y133_SLICE_X4Y133_B5Q;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C1 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C2 = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C3 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B1 = CLBLM_L_X8Y131_SLICE_X11Y131_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B2 = CLBLM_R_X7Y131_SLICE_X8Y131_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B3 = CLBLM_R_X5Y136_SLICE_X6Y136_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B6 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D1 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D2 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C2 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C4 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C5 = CLBLM_R_X3Y138_SLICE_X3Y138_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D4 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D5 = CLBLM_R_X11Y141_SLICE_X14Y141_BO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D6 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D2 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D3 = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D4 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D5 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D6 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A1 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A2 = CLBLM_R_X7Y138_SLICE_X8Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A3 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A4 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B1 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B5 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C1 = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C2 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C3 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C4 = CLBLM_R_X7Y140_SLICE_X9Y140_C5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C5 = CLBLM_L_X8Y138_SLICE_X11Y138_BO5;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C6 = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D2 = CLBLL_L_X4Y138_SLICE_X5Y138_C5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D3 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D5 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D6 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A2 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A4 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A5 = CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_AX = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B1 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B2 = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B3 = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B4 = CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B5 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B6 = CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_BX = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C1 = CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C2 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C4 = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C6 = CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_CX = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D1 = CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D2 = CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D4 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D6 = CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_DX = CLBLM_L_X8Y139_SLICE_X10Y139_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B5 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLM_R_X3Y139_SLICE_X2Y139_DO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D1 = CLBLM_R_X3Y129_SLICE_X3Y129_A5Q;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C3 = CLBLM_L_X8Y134_SLICE_X10Y134_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A2 = CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A3 = CLBLM_R_X7Y143_SLICE_X9Y143_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A4 = CLBLM_R_X3Y129_SLICE_X3Y129_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A6 = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B2 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B3 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B5 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B6 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C1 = CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C2 = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C3 = CLBLM_R_X5Y140_SLICE_X7Y140_DQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C5 = CLBLM_R_X3Y137_SLICE_X2Y137_DQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C6 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A4 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A5 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D1 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D2 = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D3 = CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D5 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D6 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D4 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A2 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A4 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A5 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A6 = CLBLL_L_X4Y133_SLICE_X5Y133_CQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_AX = CLBLM_L_X10Y141_SLICE_X13Y141_CO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B3 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B4 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A4 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C1 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C2 = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C3 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C5 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C6 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B4 = CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B5 = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D1 = CLBLM_R_X3Y138_SLICE_X3Y138_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D2 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D3 = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D5 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D6 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B6 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C1 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C2 = CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C3 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C5 = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X2Y137_SLICE_X0Y137_AO5;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A1 = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A3 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A4 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A5 = CLBLM_L_X8Y134_SLICE_X10Y134_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A6 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B1 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B2 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B3 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B5 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C2 = CLBLM_R_X7Y140_SLICE_X9Y140_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C3 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C5 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D1 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D3 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D2 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D3 = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D4 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D4 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D5 = CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A6 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D6 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A1 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A2 = CLBLM_L_X10Y139_SLICE_X13Y139_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A4 = CLBLM_R_X5Y137_SLICE_X6Y137_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A6 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B2 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B4 = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B5 = CLBLM_R_X11Y137_SLICE_X14Y137_A5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C1 = CLBLM_R_X7Y136_SLICE_X9Y136_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C2 = CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C3 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C4 = CLBLM_R_X3Y139_SLICE_X3Y139_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A2 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A4 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A6 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D1 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D2 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D4 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D5 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D6 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A1 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A2 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A3 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A5 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A1 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A4 = CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A5 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A6 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_AX = CLBLM_R_X7Y133_SLICE_X9Y133_CO5;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B4 = CLBLM_R_X7Y141_SLICE_X9Y141_C5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B2 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B4 = CLBLL_L_X4Y133_SLICE_X4Y133_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B5 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B5 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B6 = CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C1 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C2 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C4 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C5 = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D1 = CLBLM_R_X3Y135_SLICE_X2Y135_BQ;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_A1 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_A2 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_A3 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_A4 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_A5 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_A6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D2 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D4 = CLBLL_L_X4Y139_SLICE_X5Y139_DQ;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_B1 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_B2 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_B3 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_B4 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_B5 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_B6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A2 = CLBLM_R_X7Y134_SLICE_X8Y134_D5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A3 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_C1 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_C2 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_C3 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_C4 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_C5 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_C6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A6 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_AX = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B2 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C4 = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B3 = CLBLM_R_X3Y133_SLICE_X3Y133_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B4 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C5 = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_D2 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_D1 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_D3 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_D5 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_D6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C6 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X3Y165_SLICE_X3Y165_D4 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C2 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C3 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C4 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_A1 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_A2 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_A3 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_A4 = CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_A5 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_A6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D1 = CLBLM_R_X7Y141_SLICE_X8Y141_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D2 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_B1 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_B2 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_B3 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_B4 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_B5 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_B6 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_C1 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_C2 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_C3 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_C4 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_C5 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_C6 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_D1 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_D2 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_D3 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_D4 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_D5 = 1'b1;
  assign CLBLM_R_X3Y165_SLICE_X2Y165_D6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A2 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A3 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A5 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A6 = CLBLM_R_X5Y139_SLICE_X6Y139_A5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B2 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B3 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B5 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B6 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C1 = CLBLM_R_X5Y137_SLICE_X6Y137_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C2 = CLBLM_R_X5Y140_SLICE_X6Y140_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C3 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D2 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D3 = CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D6 = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A1 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A2 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A3 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A5 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A6 = CLBLM_R_X7Y140_SLICE_X8Y140_DQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B1 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B2 = CLBLM_R_X3Y134_SLICE_X2Y134_DQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B3 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B5 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C2 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C3 = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C5 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D1 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D3 = CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D4 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D6 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLL_L_X2Y139_SLICE_X0Y139_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A2 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A3 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A5 = CLBLM_R_X5Y135_SLICE_X7Y135_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B1 = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B2 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B3 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B5 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B6 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C1 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C2 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C3 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C5 = CLBLL_L_X4Y137_SLICE_X5Y137_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D1 = CLBLM_R_X5Y134_SLICE_X7Y134_C5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D2 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D3 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D5 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A1 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A3 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A6 = CLBLM_R_X5Y132_SLICE_X6Y132_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B1 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B2 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B3 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B5 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B6 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C2 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C3 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C4 = CLBLM_R_X7Y134_SLICE_X9Y134_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C5 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C6 = CLBLM_R_X7Y134_SLICE_X8Y134_D5Q;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y138_SLICE_X3Y138_B5Q;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = CLBLM_R_X5Y141_SLICE_X6Y141_C5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D2 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D3 = CLBLM_R_X5Y140_SLICE_X6Y140_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D4 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D5 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = CLBLL_L_X2Y135_SLICE_X1Y135_CQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A5 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A6 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_AX = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D1 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D2 = CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B1 = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D3 = CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B2 = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D4 = CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B3 = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D5 = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B4 = CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C2 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D6 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C3 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B5 = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B6 = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A1 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A2 = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A5 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A6 = CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B1 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B2 = CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B3 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B4 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B5 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B6 = CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C1 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C2 = CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C3 = CLBLM_R_X5Y144_SLICE_X7Y144_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C4 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C5 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C6 = CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D2 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D4 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A1 = CLBLM_R_X3Y136_SLICE_X3Y136_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A2 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A5 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A6 = CLBLM_R_X7Y141_SLICE_X9Y141_DQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B2 = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B4 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B5 = CLBLM_R_X5Y142_SLICE_X7Y142_DQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D2 = CLBLL_L_X4Y139_SLICE_X5Y139_DQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C2 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C3 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C4 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C6 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D6 = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D1 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D2 = CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D4 = CLBLM_R_X5Y138_SLICE_X7Y138_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D5 = CLBLM_R_X5Y138_SLICE_X7Y138_B5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A1 = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A2 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A3 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A5 = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A6 = 1'b1;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B2 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B3 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B5 = CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B6 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D4 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D5 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_BX = CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C1 = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C2 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C3 = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C6 = CLBLM_R_X7Y134_SLICE_X8Y134_DQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D2 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D3 = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D4 = CLBLM_L_X8Y138_SLICE_X11Y138_BO5;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D5 = CLBLL_L_X4Y135_SLICE_X4Y135_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D6 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A1 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A3 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A4 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A5 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A6 = CLBLM_R_X7Y140_SLICE_X9Y140_C5Q;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X2Y139_SLICE_X0Y139_BQ;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y138_SLICE_X5Y138_CQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_AX = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B1 = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B2 = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B3 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B4 = CLBLM_R_X5Y133_SLICE_X7Y133_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B5 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B6 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_BX = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C1 = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C2 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C3 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C4 = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C5 = CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C6 = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D1 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D3 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D4 = CLBLM_R_X5Y140_SLICE_X6Y140_C5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D5 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D6 = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C4 = CLBLM_R_X11Y140_SLICE_X14Y140_BO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C4 = CLBLM_R_X7Y129_SLICE_X9Y129_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C5 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C5 = CLBLM_R_X5Y137_SLICE_X6Y137_B5Q;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D2 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C6 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A1 = CLBLM_R_X5Y144_SLICE_X7Y144_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A2 = CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A3 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A4 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A5 = CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D2 = CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B5 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A1 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A3 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A4 = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A6 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D6 = CLBLM_R_X3Y135_SLICE_X2Y135_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B1 = CLBLL_L_X4Y140_SLICE_X5Y140_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B2 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B3 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B4 = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B5 = CLBLL_L_X2Y137_SLICE_X0Y137_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C1 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C2 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C3 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C3 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D4 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D6 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C5 = CLBLL_L_X2Y139_SLICE_X0Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A1 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A3 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A6 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B1 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B2 = CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_DQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B5 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C1 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C2 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C3 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C5 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D5 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D1 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D2 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D3 = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D4 = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D6 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A1 = CLBLM_R_X7Y136_SLICE_X8Y136_B5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A3 = CLBLM_R_X5Y135_SLICE_X6Y135_CQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A4 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A5 = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B1 = CLBLL_L_X4Y131_SLICE_X5Y131_D5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B2 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B3 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B5 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B6 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C1 = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C2 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C3 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C4 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C5 = CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C6 = CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B2 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D1 = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D2 = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D3 = CLBLM_R_X3Y134_SLICE_X2Y134_DQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D5 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B3 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D6 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D2 = CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A1 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A2 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A2 = CLBLM_L_X8Y140_SLICE_X11Y140_DQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A3 = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A3 = CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A4 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A6 = CLBLL_L_X2Y135_SLICE_X1Y135_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A4 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B2 = CLBLL_L_X2Y138_SLICE_X1Y138_BQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B3 = CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B4 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B5 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D5 = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B3 = CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B6 = CLBLL_L_X2Y135_SLICE_X1Y135_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B6 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C1 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C2 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C4 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C5 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C3 = CLBLL_L_X2Y135_SLICE_X1Y135_BQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C5 = CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C6 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D6 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D4 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D3 = CLBLL_L_X2Y135_SLICE_X1Y135_DQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D4 = CLBLM_R_X3Y134_SLICE_X3Y134_DQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D5 = CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A5 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A6 = CLBLM_R_X7Y141_SLICE_X9Y141_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A2 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B1 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B2 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B3 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B4 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B5 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D4 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X11Y139_SLICE_X14Y139_CO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C1 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C3 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C4 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D6 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D4 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D6 = CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A1 = CLBLL_L_X4Y136_SLICE_X5Y136_B5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A2 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A4 = CLBLM_R_X3Y129_SLICE_X3Y129_A5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A5 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B1 = CLBLM_R_X7Y140_SLICE_X9Y140_DQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B2 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B3 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B5 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B6 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D6 = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C1 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C2 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C3 = CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C4 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C6 = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D2 = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D3 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D4 = CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D5 = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D6 = CLBLM_R_X3Y137_SLICE_X2Y137_D5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A6 = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A2 = CLBLM_R_X5Y135_SLICE_X6Y135_C5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A3 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A4 = CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A5 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A6 = CLBLL_L_X4Y131_SLICE_X5Y131_DQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B1 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B2 = CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B3 = CLBLM_R_X5Y136_SLICE_X7Y136_C5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B5 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C1 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C2 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C3 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B1 = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_DQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B2 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y197_IOB_X0Y198_O = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B3 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D2 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D4 = CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D5 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D6 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B5 = CLBLM_L_X8Y132_SLICE_X10Y132_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B6 = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C1 = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C2 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B4 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C3 = CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C5 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C6 = CLBLM_L_X10Y140_SLICE_X12Y140_DO5;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D2 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D5 = CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A1 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A2 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A3 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A5 = CLBLM_R_X5Y135_SLICE_X6Y135_CQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A6 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B1 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B2 = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B4 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B5 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C1 = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C2 = CLBLM_R_X5Y135_SLICE_X6Y135_DQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C3 = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C4 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C5 = CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B5 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C6 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B6 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D1 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D2 = CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D3 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D4 = CLBLM_L_X10Y137_SLICE_X12Y137_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D5 = CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D6 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A1 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A2 = CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A3 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A4 = CLBLM_R_X3Y138_SLICE_X3Y138_D5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B1 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B2 = CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B3 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B5 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C1 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C2 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C3 = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C4 = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C5 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C4 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C6 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C5 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_C5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D2 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D3 = CLBLL_L_X4Y139_SLICE_X5Y139_D5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A1 = CLBLM_R_X3Y138_SLICE_X2Y138_DQ;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A2 = CLBLM_R_X3Y137_SLICE_X2Y137_D5Q;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A3 = CLBLL_L_X2Y137_SLICE_X0Y137_AQ;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A5 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D5 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D6 = CLBLM_R_X3Y138_SLICE_X3Y138_D5Q;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B1 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B2 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B3 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B4 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B5 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B6 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C1 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C2 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C3 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C4 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C5 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C6 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D1 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D2 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D3 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D4 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D5 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D6 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A1 = CLBLM_R_X3Y134_SLICE_X3Y134_DQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A2 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A3 = CLBLL_L_X2Y137_SLICE_X1Y137_AQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A4 = CLBLL_L_X2Y137_SLICE_X1Y137_CQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = CLBLM_R_X3Y133_SLICE_X2Y133_DO5;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B1 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B2 = CLBLL_L_X2Y137_SLICE_X1Y137_BQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B3 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B5 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B6 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C1 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C2 = CLBLL_L_X2Y137_SLICE_X1Y137_CQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C4 = CLBLM_R_X5Y136_SLICE_X7Y136_A5Q;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C6 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D1 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D2 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D3 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D4 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D5 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D6 = 1'b1;
endmodule
